module BoothEncoder_radix4( // @[:@3.2]
  output [2:0]  io_eB_0, // @[:@6.4]
  output [2:0]  io_eB_1, // @[:@6.4]
  output [2:0]  io_eB_2, // @[:@6.4]
  output [2:0]  io_eB_3, // @[:@6.4]
  output [2:0]  io_eB_4, // @[:@6.4]
  output [2:0]  io_eB_5, // @[:@6.4]
  output [2:0]  io_eB_6, // @[:@6.4]
  output [2:0]  io_eB_7, // @[:@6.4]
  input  [15:0] io_B // @[:@6.4]
);
  wire  _T_33; // @[RA_Mul.scala 35:28:@8.4]
  wire  _T_34; // @[RA_Mul.scala 35:28:@9.4]
  wire  _T_35; // @[RA_Mul.scala 35:28:@10.4]
  wire  _T_36; // @[RA_Mul.scala 35:28:@11.4]
  wire  _T_37; // @[RA_Mul.scala 35:28:@12.4]
  wire  _T_38; // @[RA_Mul.scala 35:28:@13.4]
  wire  _T_39; // @[RA_Mul.scala 35:28:@14.4]
  wire  _T_40; // @[RA_Mul.scala 35:28:@15.4]
  wire  _T_41; // @[RA_Mul.scala 35:28:@16.4]
  wire  _T_42; // @[RA_Mul.scala 35:28:@17.4]
  wire  _T_43; // @[RA_Mul.scala 35:28:@18.4]
  wire  _T_44; // @[RA_Mul.scala 35:28:@19.4]
  wire  _T_45; // @[RA_Mul.scala 35:28:@20.4]
  wire  _T_46; // @[RA_Mul.scala 35:28:@21.4]
  wire  _T_47; // @[RA_Mul.scala 35:28:@22.4]
  wire  _T_48; // @[RA_Mul.scala 35:28:@23.4]
  wire [1:0] _T_74; // @[RA_Mul.scala 35:51:@42.4]
  wire [1:0] _T_75; // @[RA_Mul.scala 35:51:@43.4]
  wire [3:0] _T_76; // @[RA_Mul.scala 35:51:@44.4]
  wire [1:0] _T_77; // @[RA_Mul.scala 35:51:@45.4]
  wire [1:0] _T_78; // @[RA_Mul.scala 35:51:@46.4]
  wire [3:0] _T_79; // @[RA_Mul.scala 35:51:@47.4]
  wire [7:0] _T_80; // @[RA_Mul.scala 35:51:@48.4]
  wire [1:0] _T_81; // @[RA_Mul.scala 35:51:@49.4]
  wire [1:0] _T_82; // @[RA_Mul.scala 35:51:@50.4]
  wire [3:0] _T_83; // @[RA_Mul.scala 35:51:@51.4]
  wire [1:0] _T_84; // @[RA_Mul.scala 35:51:@52.4]
  wire [1:0] _T_85; // @[RA_Mul.scala 35:51:@53.4]
  wire [2:0] _T_86; // @[RA_Mul.scala 35:51:@54.4]
  wire [4:0] _T_87; // @[RA_Mul.scala 35:51:@55.4]
  wire [8:0] _T_88; // @[RA_Mul.scala 35:51:@56.4]
  wire [16:0] B_ext; // @[RA_Mul.scala 35:51:@57.4]
  wire  _T_98; // @[RA_Mul.scala 39:24:@59.4]
  wire  _T_99; // @[RA_Mul.scala 39:37:@60.4]
  wire  _T_100; // @[RA_Mul.scala 39:30:@61.4]
  wire  _T_101; // @[RA_Mul.scala 40:25:@63.4]
  wire  _T_103; // @[RA_Mul.scala 40:36:@65.4]
  wire  _T_104; // @[RA_Mul.scala 40:33:@66.4]
  wire  _T_106; // @[RA_Mul.scala 40:54:@68.4]
  wire  _T_107; // @[RA_Mul.scala 40:51:@69.4]
  wire  _T_109; // @[RA_Mul.scala 40:70:@71.4]
  wire  _T_111; // @[RA_Mul.scala 40:85:@73.4]
  wire  _T_113; // @[RA_Mul.scala 40:100:@75.4]
  wire  _T_114; // @[RA_Mul.scala 40:66:@76.4]
  wire [1:0] _T_116; // @[RA_Mul.scala 42:25:@80.4]
  wire  _T_129; // @[RA_Mul.scala 39:30:@86.4]
  wire  _T_130; // @[RA_Mul.scala 40:25:@88.4]
  wire  _T_133; // @[RA_Mul.scala 40:33:@91.4]
  wire  _T_136; // @[RA_Mul.scala 40:51:@94.4]
  wire  _T_138; // @[RA_Mul.scala 40:70:@96.4]
  wire  _T_140; // @[RA_Mul.scala 40:85:@98.4]
  wire  _T_142; // @[RA_Mul.scala 40:100:@100.4]
  wire  _T_143; // @[RA_Mul.scala 40:66:@101.4]
  wire [1:0] _T_145; // @[RA_Mul.scala 42:25:@105.4]
  wire  _T_158; // @[RA_Mul.scala 39:30:@111.4]
  wire  _T_159; // @[RA_Mul.scala 40:25:@113.4]
  wire  _T_162; // @[RA_Mul.scala 40:33:@116.4]
  wire  _T_165; // @[RA_Mul.scala 40:51:@119.4]
  wire  _T_167; // @[RA_Mul.scala 40:70:@121.4]
  wire  _T_169; // @[RA_Mul.scala 40:85:@123.4]
  wire  _T_171; // @[RA_Mul.scala 40:100:@125.4]
  wire  _T_172; // @[RA_Mul.scala 40:66:@126.4]
  wire [1:0] _T_174; // @[RA_Mul.scala 42:25:@130.4]
  wire  _T_187; // @[RA_Mul.scala 39:30:@136.4]
  wire  _T_188; // @[RA_Mul.scala 40:25:@138.4]
  wire  _T_191; // @[RA_Mul.scala 40:33:@141.4]
  wire  _T_194; // @[RA_Mul.scala 40:51:@144.4]
  wire  _T_196; // @[RA_Mul.scala 40:70:@146.4]
  wire  _T_198; // @[RA_Mul.scala 40:85:@148.4]
  wire  _T_200; // @[RA_Mul.scala 40:100:@150.4]
  wire  _T_201; // @[RA_Mul.scala 40:66:@151.4]
  wire [1:0] _T_203; // @[RA_Mul.scala 42:25:@155.4]
  wire  _T_216; // @[RA_Mul.scala 39:30:@161.4]
  wire  _T_217; // @[RA_Mul.scala 40:25:@163.4]
  wire  _T_220; // @[RA_Mul.scala 40:33:@166.4]
  wire  _T_223; // @[RA_Mul.scala 40:51:@169.4]
  wire  _T_225; // @[RA_Mul.scala 40:70:@171.4]
  wire  _T_227; // @[RA_Mul.scala 40:85:@173.4]
  wire  _T_229; // @[RA_Mul.scala 40:100:@175.4]
  wire  _T_230; // @[RA_Mul.scala 40:66:@176.4]
  wire [1:0] _T_232; // @[RA_Mul.scala 42:25:@180.4]
  wire  _T_245; // @[RA_Mul.scala 39:30:@186.4]
  wire  _T_246; // @[RA_Mul.scala 40:25:@188.4]
  wire  _T_249; // @[RA_Mul.scala 40:33:@191.4]
  wire  _T_252; // @[RA_Mul.scala 40:51:@194.4]
  wire  _T_254; // @[RA_Mul.scala 40:70:@196.4]
  wire  _T_256; // @[RA_Mul.scala 40:85:@198.4]
  wire  _T_258; // @[RA_Mul.scala 40:100:@200.4]
  wire  _T_259; // @[RA_Mul.scala 40:66:@201.4]
  wire [1:0] _T_261; // @[RA_Mul.scala 42:25:@205.4]
  wire  _T_274; // @[RA_Mul.scala 39:30:@211.4]
  wire  _T_275; // @[RA_Mul.scala 40:25:@213.4]
  wire  _T_278; // @[RA_Mul.scala 40:33:@216.4]
  wire  _T_281; // @[RA_Mul.scala 40:51:@219.4]
  wire  _T_283; // @[RA_Mul.scala 40:70:@221.4]
  wire  _T_285; // @[RA_Mul.scala 40:85:@223.4]
  wire  _T_287; // @[RA_Mul.scala 40:100:@225.4]
  wire  _T_288; // @[RA_Mul.scala 40:66:@226.4]
  wire [1:0] _T_290; // @[RA_Mul.scala 42:25:@230.4]
  wire  _T_303; // @[RA_Mul.scala 39:30:@236.4]
  wire  _T_304; // @[RA_Mul.scala 40:25:@238.4]
  wire  _T_307; // @[RA_Mul.scala 40:33:@241.4]
  wire  _T_310; // @[RA_Mul.scala 40:51:@244.4]
  wire  _T_312; // @[RA_Mul.scala 40:70:@246.4]
  wire  _T_314; // @[RA_Mul.scala 40:85:@248.4]
  wire  _T_316; // @[RA_Mul.scala 40:100:@250.4]
  wire  _T_317; // @[RA_Mul.scala 40:66:@251.4]
  wire [1:0] _T_319; // @[RA_Mul.scala 42:25:@255.4]
  assign _T_33 = io_B[0]; // @[RA_Mul.scala 35:28:@8.4]
  assign _T_34 = io_B[1]; // @[RA_Mul.scala 35:28:@9.4]
  assign _T_35 = io_B[2]; // @[RA_Mul.scala 35:28:@10.4]
  assign _T_36 = io_B[3]; // @[RA_Mul.scala 35:28:@11.4]
  assign _T_37 = io_B[4]; // @[RA_Mul.scala 35:28:@12.4]
  assign _T_38 = io_B[5]; // @[RA_Mul.scala 35:28:@13.4]
  assign _T_39 = io_B[6]; // @[RA_Mul.scala 35:28:@14.4]
  assign _T_40 = io_B[7]; // @[RA_Mul.scala 35:28:@15.4]
  assign _T_41 = io_B[8]; // @[RA_Mul.scala 35:28:@16.4]
  assign _T_42 = io_B[9]; // @[RA_Mul.scala 35:28:@17.4]
  assign _T_43 = io_B[10]; // @[RA_Mul.scala 35:28:@18.4]
  assign _T_44 = io_B[11]; // @[RA_Mul.scala 35:28:@19.4]
  assign _T_45 = io_B[12]; // @[RA_Mul.scala 35:28:@20.4]
  assign _T_46 = io_B[13]; // @[RA_Mul.scala 35:28:@21.4]
  assign _T_47 = io_B[14]; // @[RA_Mul.scala 35:28:@22.4]
  assign _T_48 = io_B[15]; // @[RA_Mul.scala 35:28:@23.4]
  assign _T_74 = {_T_34,_T_33}; // @[RA_Mul.scala 35:51:@42.4]
  assign _T_75 = {_T_36,_T_35}; // @[RA_Mul.scala 35:51:@43.4]
  assign _T_76 = {_T_75,_T_74}; // @[RA_Mul.scala 35:51:@44.4]
  assign _T_77 = {_T_38,_T_37}; // @[RA_Mul.scala 35:51:@45.4]
  assign _T_78 = {_T_40,_T_39}; // @[RA_Mul.scala 35:51:@46.4]
  assign _T_79 = {_T_78,_T_77}; // @[RA_Mul.scala 35:51:@47.4]
  assign _T_80 = {_T_79,_T_76}; // @[RA_Mul.scala 35:51:@48.4]
  assign _T_81 = {_T_42,_T_41}; // @[RA_Mul.scala 35:51:@49.4]
  assign _T_82 = {_T_44,_T_43}; // @[RA_Mul.scala 35:51:@50.4]
  assign _T_83 = {_T_82,_T_81}; // @[RA_Mul.scala 35:51:@51.4]
  assign _T_84 = {_T_46,_T_45}; // @[RA_Mul.scala 35:51:@52.4]
  assign _T_85 = {1'h0,_T_48}; // @[RA_Mul.scala 35:51:@53.4]
  assign _T_86 = {_T_85,_T_47}; // @[RA_Mul.scala 35:51:@54.4]
  assign _T_87 = {_T_86,_T_84}; // @[RA_Mul.scala 35:51:@55.4]
  assign _T_88 = {_T_87,_T_83}; // @[RA_Mul.scala 35:51:@56.4]
  assign B_ext = {_T_88,_T_80}; // @[RA_Mul.scala 35:51:@57.4]
  assign _T_98 = B_ext[1]; // @[RA_Mul.scala 39:24:@59.4]
  assign _T_99 = B_ext[0]; // @[RA_Mul.scala 39:37:@60.4]
  assign _T_100 = _T_98 ^ _T_99; // @[RA_Mul.scala 39:30:@61.4]
  assign _T_101 = B_ext[2]; // @[RA_Mul.scala 40:25:@63.4]
  assign _T_103 = ~ _T_98; // @[RA_Mul.scala 40:36:@65.4]
  assign _T_104 = _T_101 & _T_103; // @[RA_Mul.scala 40:33:@66.4]
  assign _T_106 = ~ _T_99; // @[RA_Mul.scala 40:54:@68.4]
  assign _T_107 = _T_104 & _T_106; // @[RA_Mul.scala 40:51:@69.4]
  assign _T_109 = ~ _T_101; // @[RA_Mul.scala 40:70:@71.4]
  assign _T_111 = _T_109 & _T_98; // @[RA_Mul.scala 40:85:@73.4]
  assign _T_113 = _T_111 & _T_99; // @[RA_Mul.scala 40:100:@75.4]
  assign _T_114 = _T_107 | _T_113; // @[RA_Mul.scala 40:66:@76.4]
  assign _T_116 = {_T_101,_T_114}; // @[RA_Mul.scala 42:25:@80.4]
  assign _T_129 = _T_101 ^ _T_98; // @[RA_Mul.scala 39:30:@86.4]
  assign _T_130 = B_ext[3]; // @[RA_Mul.scala 40:25:@88.4]
  assign _T_133 = _T_130 & _T_109; // @[RA_Mul.scala 40:33:@91.4]
  assign _T_136 = _T_133 & _T_103; // @[RA_Mul.scala 40:51:@94.4]
  assign _T_138 = ~ _T_130; // @[RA_Mul.scala 40:70:@96.4]
  assign _T_140 = _T_138 & _T_101; // @[RA_Mul.scala 40:85:@98.4]
  assign _T_142 = _T_140 & _T_98; // @[RA_Mul.scala 40:100:@100.4]
  assign _T_143 = _T_136 | _T_142; // @[RA_Mul.scala 40:66:@101.4]
  assign _T_145 = {_T_130,_T_143}; // @[RA_Mul.scala 42:25:@105.4]
  assign _T_158 = _T_130 ^ _T_101; // @[RA_Mul.scala 39:30:@111.4]
  assign _T_159 = B_ext[4]; // @[RA_Mul.scala 40:25:@113.4]
  assign _T_162 = _T_159 & _T_138; // @[RA_Mul.scala 40:33:@116.4]
  assign _T_165 = _T_162 & _T_109; // @[RA_Mul.scala 40:51:@119.4]
  assign _T_167 = ~ _T_159; // @[RA_Mul.scala 40:70:@121.4]
  assign _T_169 = _T_167 & _T_130; // @[RA_Mul.scala 40:85:@123.4]
  assign _T_171 = _T_169 & _T_101; // @[RA_Mul.scala 40:100:@125.4]
  assign _T_172 = _T_165 | _T_171; // @[RA_Mul.scala 40:66:@126.4]
  assign _T_174 = {_T_159,_T_172}; // @[RA_Mul.scala 42:25:@130.4]
  assign _T_187 = _T_159 ^ _T_130; // @[RA_Mul.scala 39:30:@136.4]
  assign _T_188 = B_ext[5]; // @[RA_Mul.scala 40:25:@138.4]
  assign _T_191 = _T_188 & _T_167; // @[RA_Mul.scala 40:33:@141.4]
  assign _T_194 = _T_191 & _T_138; // @[RA_Mul.scala 40:51:@144.4]
  assign _T_196 = ~ _T_188; // @[RA_Mul.scala 40:70:@146.4]
  assign _T_198 = _T_196 & _T_159; // @[RA_Mul.scala 40:85:@148.4]
  assign _T_200 = _T_198 & _T_130; // @[RA_Mul.scala 40:100:@150.4]
  assign _T_201 = _T_194 | _T_200; // @[RA_Mul.scala 40:66:@151.4]
  assign _T_203 = {_T_188,_T_201}; // @[RA_Mul.scala 42:25:@155.4]
  assign _T_216 = _T_188 ^ _T_159; // @[RA_Mul.scala 39:30:@161.4]
  assign _T_217 = B_ext[6]; // @[RA_Mul.scala 40:25:@163.4]
  assign _T_220 = _T_217 & _T_196; // @[RA_Mul.scala 40:33:@166.4]
  assign _T_223 = _T_220 & _T_167; // @[RA_Mul.scala 40:51:@169.4]
  assign _T_225 = ~ _T_217; // @[RA_Mul.scala 40:70:@171.4]
  assign _T_227 = _T_225 & _T_188; // @[RA_Mul.scala 40:85:@173.4]
  assign _T_229 = _T_227 & _T_159; // @[RA_Mul.scala 40:100:@175.4]
  assign _T_230 = _T_223 | _T_229; // @[RA_Mul.scala 40:66:@176.4]
  assign _T_232 = {_T_217,_T_230}; // @[RA_Mul.scala 42:25:@180.4]
  assign _T_245 = _T_217 ^ _T_188; // @[RA_Mul.scala 39:30:@186.4]
  assign _T_246 = B_ext[7]; // @[RA_Mul.scala 40:25:@188.4]
  assign _T_249 = _T_246 & _T_225; // @[RA_Mul.scala 40:33:@191.4]
  assign _T_252 = _T_249 & _T_196; // @[RA_Mul.scala 40:51:@194.4]
  assign _T_254 = ~ _T_246; // @[RA_Mul.scala 40:70:@196.4]
  assign _T_256 = _T_254 & _T_217; // @[RA_Mul.scala 40:85:@198.4]
  assign _T_258 = _T_256 & _T_188; // @[RA_Mul.scala 40:100:@200.4]
  assign _T_259 = _T_252 | _T_258; // @[RA_Mul.scala 40:66:@201.4]
  assign _T_261 = {_T_246,_T_259}; // @[RA_Mul.scala 42:25:@205.4]
  assign _T_274 = _T_246 ^ _T_217; // @[RA_Mul.scala 39:30:@211.4]
  assign _T_275 = B_ext[8]; // @[RA_Mul.scala 40:25:@213.4]
  assign _T_278 = _T_275 & _T_254; // @[RA_Mul.scala 40:33:@216.4]
  assign _T_281 = _T_278 & _T_225; // @[RA_Mul.scala 40:51:@219.4]
  assign _T_283 = ~ _T_275; // @[RA_Mul.scala 40:70:@221.4]
  assign _T_285 = _T_283 & _T_246; // @[RA_Mul.scala 40:85:@223.4]
  assign _T_287 = _T_285 & _T_217; // @[RA_Mul.scala 40:100:@225.4]
  assign _T_288 = _T_281 | _T_287; // @[RA_Mul.scala 40:66:@226.4]
  assign _T_290 = {_T_275,_T_288}; // @[RA_Mul.scala 42:25:@230.4]
  assign _T_303 = _T_275 ^ _T_246; // @[RA_Mul.scala 39:30:@236.4]
  assign _T_304 = B_ext[9]; // @[RA_Mul.scala 40:25:@238.4]
  assign _T_307 = _T_304 & _T_283; // @[RA_Mul.scala 40:33:@241.4]
  assign _T_310 = _T_307 & _T_254; // @[RA_Mul.scala 40:51:@244.4]
  assign _T_312 = ~ _T_304; // @[RA_Mul.scala 40:70:@246.4]
  assign _T_314 = _T_312 & _T_275; // @[RA_Mul.scala 40:85:@248.4]
  assign _T_316 = _T_314 & _T_246; // @[RA_Mul.scala 40:100:@250.4]
  assign _T_317 = _T_310 | _T_316; // @[RA_Mul.scala 40:66:@251.4]
  assign _T_319 = {_T_304,_T_317}; // @[RA_Mul.scala 42:25:@255.4]
  assign io_eB_0 = {_T_116,_T_100}; // @[RA_Mul.scala 42:15:@82.4]
  assign io_eB_1 = {_T_145,_T_129}; // @[RA_Mul.scala 42:15:@107.4]
  assign io_eB_2 = {_T_174,_T_158}; // @[RA_Mul.scala 42:15:@132.4]
  assign io_eB_3 = {_T_203,_T_187}; // @[RA_Mul.scala 42:15:@157.4]
  assign io_eB_4 = {_T_232,_T_216}; // @[RA_Mul.scala 42:15:@182.4]
  assign io_eB_5 = {_T_261,_T_245}; // @[RA_Mul.scala 42:15:@207.4]
  assign io_eB_6 = {_T_290,_T_274}; // @[RA_Mul.scala 42:15:@232.4]
  assign io_eB_7 = {_T_319,_T_303}; // @[RA_Mul.scala 42:15:@257.4]
endmodule
module PPGen( // @[:@259.2]
  output [15:0] io_PP_0, // @[:@262.4]
  output [15:0] io_PP_1, // @[:@262.4]
  output [15:0] io_PP_2, // @[:@262.4]
  output [15:0] io_PP_3, // @[:@262.4]
  output [15:0] io_PP_4, // @[:@262.4]
  output [15:0] io_PP_5, // @[:@262.4]
  output [15:0] io_PP_6, // @[:@262.4]
  output [15:0] io_PP_7, // @[:@262.4]
  output [7:0]  io_SC, // @[:@262.4]
  output [7:0]  io_S, // @[:@262.4]
  input  [2:0]  io_eB_0, // @[:@262.4]
  input  [2:0]  io_eB_1, // @[:@262.4]
  input  [2:0]  io_eB_2, // @[:@262.4]
  input  [2:0]  io_eB_3, // @[:@262.4]
  input  [2:0]  io_eB_4, // @[:@262.4]
  input  [2:0]  io_eB_5, // @[:@262.4]
  input  [2:0]  io_eB_6, // @[:@262.4]
  input  [2:0]  io_eB_7, // @[:@262.4]
  input  [15:0] io_A // @[:@262.4]
);
  wire  _T_93; // @[RA_Mul.scala 62:19:@267.4]
  wire  _T_95; // @[RA_Mul.scala 62:44:@268.4]
  wire  _T_96; // @[RA_Mul.scala 62:32:@269.4]
  wire  _T_99; // @[RA_Mul.scala 64:25:@274.6]
  wire  _T_101; // @[RA_Mul.scala 66:25:@279.8]
  wire [16:0] _GEN_40; // @[RA_Mul.scala 67:25:@281.10]
  wire [16:0] _T_102; // @[RA_Mul.scala 67:25:@281.10]
  wire [15:0] _T_103; // @[RA_Mul.scala 67:30:@282.10]
  wire  _T_105; // @[RA_Mul.scala 68:25:@286.10]
  wire [15:0] _T_106; // @[RA_Mul.scala 69:19:@288.12]
  wire  _T_108; // @[RA_Mul.scala 70:25:@292.12]
  wire [15:0] _T_111; // @[RA_Mul.scala 71:19:@296.14]
  wire [15:0] _GEN_0; // @[RA_Mul.scala 70:38:@293.12]
  wire [15:0] _GEN_1; // @[RA_Mul.scala 68:39:@287.10]
  wire [15:0] _GEN_2; // @[RA_Mul.scala 66:39:@280.8]
  wire [15:0] _GEN_3; // @[RA_Mul.scala 64:39:@275.6]
  wire  S_v_0; // @[RA_Mul.scala 76:23:@302.4]
  wire  _T_115; // @[RA_Mul.scala 77:36:@305.4]
  wire  _T_116; // @[RA_Mul.scala 77:30:@306.4]
  wire  SC_v_0; // @[RA_Mul.scala 77:16:@307.4]
  wire  _T_119; // @[RA_Mul.scala 62:19:@309.4]
  wire  _T_121; // @[RA_Mul.scala 62:44:@310.4]
  wire  _T_122; // @[RA_Mul.scala 62:32:@311.4]
  wire  _T_125; // @[RA_Mul.scala 64:25:@316.6]
  wire  _T_127; // @[RA_Mul.scala 66:25:@321.8]
  wire  _T_131; // @[RA_Mul.scala 68:25:@328.10]
  wire  _T_134; // @[RA_Mul.scala 70:25:@334.12]
  wire [15:0] _GEN_5; // @[RA_Mul.scala 70:38:@335.12]
  wire [15:0] _GEN_6; // @[RA_Mul.scala 68:39:@329.10]
  wire [15:0] _GEN_7; // @[RA_Mul.scala 66:39:@322.8]
  wire [15:0] _GEN_8; // @[RA_Mul.scala 64:39:@317.6]
  wire  S_v_1; // @[RA_Mul.scala 76:23:@344.4]
  wire  _T_142; // @[RA_Mul.scala 77:30:@348.4]
  wire  SC_v_1; // @[RA_Mul.scala 77:16:@349.4]
  wire  _T_145; // @[RA_Mul.scala 62:19:@351.4]
  wire  _T_147; // @[RA_Mul.scala 62:44:@352.4]
  wire  _T_148; // @[RA_Mul.scala 62:32:@353.4]
  wire  _T_151; // @[RA_Mul.scala 64:25:@358.6]
  wire  _T_153; // @[RA_Mul.scala 66:25:@363.8]
  wire  _T_157; // @[RA_Mul.scala 68:25:@370.10]
  wire  _T_160; // @[RA_Mul.scala 70:25:@376.12]
  wire [15:0] _GEN_10; // @[RA_Mul.scala 70:38:@377.12]
  wire [15:0] _GEN_11; // @[RA_Mul.scala 68:39:@371.10]
  wire [15:0] _GEN_12; // @[RA_Mul.scala 66:39:@364.8]
  wire [15:0] _GEN_13; // @[RA_Mul.scala 64:39:@359.6]
  wire  S_v_2; // @[RA_Mul.scala 76:23:@386.4]
  wire  _T_168; // @[RA_Mul.scala 77:30:@390.4]
  wire  SC_v_2; // @[RA_Mul.scala 77:16:@391.4]
  wire  _T_171; // @[RA_Mul.scala 62:19:@393.4]
  wire  _T_173; // @[RA_Mul.scala 62:44:@394.4]
  wire  _T_174; // @[RA_Mul.scala 62:32:@395.4]
  wire  _T_177; // @[RA_Mul.scala 64:25:@400.6]
  wire  _T_179; // @[RA_Mul.scala 66:25:@405.8]
  wire  _T_183; // @[RA_Mul.scala 68:25:@412.10]
  wire  _T_186; // @[RA_Mul.scala 70:25:@418.12]
  wire [15:0] _GEN_15; // @[RA_Mul.scala 70:38:@419.12]
  wire [15:0] _GEN_16; // @[RA_Mul.scala 68:39:@413.10]
  wire [15:0] _GEN_17; // @[RA_Mul.scala 66:39:@406.8]
  wire [15:0] _GEN_18; // @[RA_Mul.scala 64:39:@401.6]
  wire  S_v_3; // @[RA_Mul.scala 76:23:@428.4]
  wire  _T_194; // @[RA_Mul.scala 77:30:@432.4]
  wire  SC_v_3; // @[RA_Mul.scala 77:16:@433.4]
  wire  _T_197; // @[RA_Mul.scala 62:19:@435.4]
  wire  _T_199; // @[RA_Mul.scala 62:44:@436.4]
  wire  _T_200; // @[RA_Mul.scala 62:32:@437.4]
  wire  _T_203; // @[RA_Mul.scala 64:25:@442.6]
  wire  _T_205; // @[RA_Mul.scala 66:25:@447.8]
  wire  _T_209; // @[RA_Mul.scala 68:25:@454.10]
  wire  _T_212; // @[RA_Mul.scala 70:25:@460.12]
  wire [15:0] _GEN_20; // @[RA_Mul.scala 70:38:@461.12]
  wire [15:0] _GEN_21; // @[RA_Mul.scala 68:39:@455.10]
  wire [15:0] _GEN_22; // @[RA_Mul.scala 66:39:@448.8]
  wire [15:0] _GEN_23; // @[RA_Mul.scala 64:39:@443.6]
  wire  S_v_4; // @[RA_Mul.scala 76:23:@470.4]
  wire  _T_220; // @[RA_Mul.scala 77:30:@474.4]
  wire  SC_v_4; // @[RA_Mul.scala 77:16:@475.4]
  wire  _T_223; // @[RA_Mul.scala 62:19:@477.4]
  wire  _T_225; // @[RA_Mul.scala 62:44:@478.4]
  wire  _T_226; // @[RA_Mul.scala 62:32:@479.4]
  wire  _T_229; // @[RA_Mul.scala 64:25:@484.6]
  wire  _T_231; // @[RA_Mul.scala 66:25:@489.8]
  wire  _T_235; // @[RA_Mul.scala 68:25:@496.10]
  wire  _T_238; // @[RA_Mul.scala 70:25:@502.12]
  wire [15:0] _GEN_25; // @[RA_Mul.scala 70:38:@503.12]
  wire [15:0] _GEN_26; // @[RA_Mul.scala 68:39:@497.10]
  wire [15:0] _GEN_27; // @[RA_Mul.scala 66:39:@490.8]
  wire [15:0] _GEN_28; // @[RA_Mul.scala 64:39:@485.6]
  wire  S_v_5; // @[RA_Mul.scala 76:23:@512.4]
  wire  _T_246; // @[RA_Mul.scala 77:30:@516.4]
  wire  SC_v_5; // @[RA_Mul.scala 77:16:@517.4]
  wire  _T_249; // @[RA_Mul.scala 62:19:@519.4]
  wire  _T_251; // @[RA_Mul.scala 62:44:@520.4]
  wire  _T_252; // @[RA_Mul.scala 62:32:@521.4]
  wire  _T_255; // @[RA_Mul.scala 64:25:@526.6]
  wire  _T_257; // @[RA_Mul.scala 66:25:@531.8]
  wire  _T_261; // @[RA_Mul.scala 68:25:@538.10]
  wire  _T_264; // @[RA_Mul.scala 70:25:@544.12]
  wire [15:0] _GEN_30; // @[RA_Mul.scala 70:38:@545.12]
  wire [15:0] _GEN_31; // @[RA_Mul.scala 68:39:@539.10]
  wire [15:0] _GEN_32; // @[RA_Mul.scala 66:39:@532.8]
  wire [15:0] _GEN_33; // @[RA_Mul.scala 64:39:@527.6]
  wire  S_v_6; // @[RA_Mul.scala 76:23:@554.4]
  wire  _T_272; // @[RA_Mul.scala 77:30:@558.4]
  wire  SC_v_6; // @[RA_Mul.scala 77:16:@559.4]
  wire  _T_275; // @[RA_Mul.scala 62:19:@561.4]
  wire  _T_277; // @[RA_Mul.scala 62:44:@562.4]
  wire  _T_278; // @[RA_Mul.scala 62:32:@563.4]
  wire  _T_281; // @[RA_Mul.scala 64:25:@568.6]
  wire  _T_283; // @[RA_Mul.scala 66:25:@573.8]
  wire  _T_287; // @[RA_Mul.scala 68:25:@580.10]
  wire  _T_290; // @[RA_Mul.scala 70:25:@586.12]
  wire [15:0] _GEN_35; // @[RA_Mul.scala 70:38:@587.12]
  wire [15:0] _GEN_36; // @[RA_Mul.scala 68:39:@581.10]
  wire [15:0] _GEN_37; // @[RA_Mul.scala 66:39:@574.8]
  wire [15:0] _GEN_38; // @[RA_Mul.scala 64:39:@569.6]
  wire  S_v_7; // @[RA_Mul.scala 76:23:@596.4]
  wire  _T_298; // @[RA_Mul.scala 77:30:@600.4]
  wire  SC_v_7; // @[RA_Mul.scala 77:16:@601.4]
  wire [1:0] _T_300; // @[RA_Mul.scala 79:21:@603.4]
  wire [1:0] _T_301; // @[RA_Mul.scala 79:21:@604.4]
  wire [3:0] _T_302; // @[RA_Mul.scala 79:21:@605.4]
  wire [1:0] _T_303; // @[RA_Mul.scala 79:21:@606.4]
  wire [1:0] _T_304; // @[RA_Mul.scala 79:21:@607.4]
  wire [3:0] _T_305; // @[RA_Mul.scala 79:21:@608.4]
  wire [1:0] _T_307; // @[RA_Mul.scala 80:23:@611.4]
  wire [1:0] _T_308; // @[RA_Mul.scala 80:23:@612.4]
  wire [3:0] _T_309; // @[RA_Mul.scala 80:23:@613.4]
  wire [1:0] _T_310; // @[RA_Mul.scala 80:23:@614.4]
  wire [1:0] _T_311; // @[RA_Mul.scala 80:23:@615.4]
  wire [3:0] _T_312; // @[RA_Mul.scala 80:23:@616.4]
  assign _T_93 = io_eB_0 == 3'h0; // @[RA_Mul.scala 62:19:@267.4]
  assign _T_95 = io_eB_0 == 3'h4; // @[RA_Mul.scala 62:44:@268.4]
  assign _T_96 = _T_93 | _T_95; // @[RA_Mul.scala 62:32:@269.4]
  assign _T_99 = io_eB_0 == 3'h1; // @[RA_Mul.scala 64:25:@274.6]
  assign _T_101 = io_eB_0 == 3'h2; // @[RA_Mul.scala 66:25:@279.8]
  assign _GEN_40 = {{1'd0}, io_A}; // @[RA_Mul.scala 67:25:@281.10]
  assign _T_102 = _GEN_40 << 1; // @[RA_Mul.scala 67:25:@281.10]
  assign _T_103 = _T_102[15:0]; // @[RA_Mul.scala 67:30:@282.10]
  assign _T_105 = io_eB_0 == 3'h5; // @[RA_Mul.scala 68:25:@286.10]
  assign _T_106 = ~ io_A; // @[RA_Mul.scala 69:19:@288.12]
  assign _T_108 = io_eB_0 == 3'h6; // @[RA_Mul.scala 70:25:@292.12]
  assign _T_111 = ~ _T_103; // @[RA_Mul.scala 71:19:@296.14]
  assign _GEN_0 = _T_108 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@293.12]
  assign _GEN_1 = _T_105 ? _T_106 : _GEN_0; // @[RA_Mul.scala 68:39:@287.10]
  assign _GEN_2 = _T_101 ? _T_103 : _GEN_1; // @[RA_Mul.scala 66:39:@280.8]
  assign _GEN_3 = _T_99 ? io_A : _GEN_2; // @[RA_Mul.scala 64:39:@275.6]
  assign S_v_0 = io_eB_0[2]; // @[RA_Mul.scala 76:23:@302.4]
  assign _T_115 = io_A[15]; // @[RA_Mul.scala 77:36:@305.4]
  assign _T_116 = S_v_0 ^ _T_115; // @[RA_Mul.scala 77:30:@306.4]
  assign SC_v_0 = ~ _T_116; // @[RA_Mul.scala 77:16:@307.4]
  assign _T_119 = io_eB_1 == 3'h0; // @[RA_Mul.scala 62:19:@309.4]
  assign _T_121 = io_eB_1 == 3'h4; // @[RA_Mul.scala 62:44:@310.4]
  assign _T_122 = _T_119 | _T_121; // @[RA_Mul.scala 62:32:@311.4]
  assign _T_125 = io_eB_1 == 3'h1; // @[RA_Mul.scala 64:25:@316.6]
  assign _T_127 = io_eB_1 == 3'h2; // @[RA_Mul.scala 66:25:@321.8]
  assign _T_131 = io_eB_1 == 3'h5; // @[RA_Mul.scala 68:25:@328.10]
  assign _T_134 = io_eB_1 == 3'h6; // @[RA_Mul.scala 70:25:@334.12]
  assign _GEN_5 = _T_134 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@335.12]
  assign _GEN_6 = _T_131 ? _T_106 : _GEN_5; // @[RA_Mul.scala 68:39:@329.10]
  assign _GEN_7 = _T_127 ? _T_103 : _GEN_6; // @[RA_Mul.scala 66:39:@322.8]
  assign _GEN_8 = _T_125 ? io_A : _GEN_7; // @[RA_Mul.scala 64:39:@317.6]
  assign S_v_1 = io_eB_1[2]; // @[RA_Mul.scala 76:23:@344.4]
  assign _T_142 = S_v_1 ^ _T_115; // @[RA_Mul.scala 77:30:@348.4]
  assign SC_v_1 = ~ _T_142; // @[RA_Mul.scala 77:16:@349.4]
  assign _T_145 = io_eB_2 == 3'h0; // @[RA_Mul.scala 62:19:@351.4]
  assign _T_147 = io_eB_2 == 3'h4; // @[RA_Mul.scala 62:44:@352.4]
  assign _T_148 = _T_145 | _T_147; // @[RA_Mul.scala 62:32:@353.4]
  assign _T_151 = io_eB_2 == 3'h1; // @[RA_Mul.scala 64:25:@358.6]
  assign _T_153 = io_eB_2 == 3'h2; // @[RA_Mul.scala 66:25:@363.8]
  assign _T_157 = io_eB_2 == 3'h5; // @[RA_Mul.scala 68:25:@370.10]
  assign _T_160 = io_eB_2 == 3'h6; // @[RA_Mul.scala 70:25:@376.12]
  assign _GEN_10 = _T_160 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@377.12]
  assign _GEN_11 = _T_157 ? _T_106 : _GEN_10; // @[RA_Mul.scala 68:39:@371.10]
  assign _GEN_12 = _T_153 ? _T_103 : _GEN_11; // @[RA_Mul.scala 66:39:@364.8]
  assign _GEN_13 = _T_151 ? io_A : _GEN_12; // @[RA_Mul.scala 64:39:@359.6]
  assign S_v_2 = io_eB_2[2]; // @[RA_Mul.scala 76:23:@386.4]
  assign _T_168 = S_v_2 ^ _T_115; // @[RA_Mul.scala 77:30:@390.4]
  assign SC_v_2 = ~ _T_168; // @[RA_Mul.scala 77:16:@391.4]
  assign _T_171 = io_eB_3 == 3'h0; // @[RA_Mul.scala 62:19:@393.4]
  assign _T_173 = io_eB_3 == 3'h4; // @[RA_Mul.scala 62:44:@394.4]
  assign _T_174 = _T_171 | _T_173; // @[RA_Mul.scala 62:32:@395.4]
  assign _T_177 = io_eB_3 == 3'h1; // @[RA_Mul.scala 64:25:@400.6]
  assign _T_179 = io_eB_3 == 3'h2; // @[RA_Mul.scala 66:25:@405.8]
  assign _T_183 = io_eB_3 == 3'h5; // @[RA_Mul.scala 68:25:@412.10]
  assign _T_186 = io_eB_3 == 3'h6; // @[RA_Mul.scala 70:25:@418.12]
  assign _GEN_15 = _T_186 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@419.12]
  assign _GEN_16 = _T_183 ? _T_106 : _GEN_15; // @[RA_Mul.scala 68:39:@413.10]
  assign _GEN_17 = _T_179 ? _T_103 : _GEN_16; // @[RA_Mul.scala 66:39:@406.8]
  assign _GEN_18 = _T_177 ? io_A : _GEN_17; // @[RA_Mul.scala 64:39:@401.6]
  assign S_v_3 = io_eB_3[2]; // @[RA_Mul.scala 76:23:@428.4]
  assign _T_194 = S_v_3 ^ _T_115; // @[RA_Mul.scala 77:30:@432.4]
  assign SC_v_3 = ~ _T_194; // @[RA_Mul.scala 77:16:@433.4]
  assign _T_197 = io_eB_4 == 3'h0; // @[RA_Mul.scala 62:19:@435.4]
  assign _T_199 = io_eB_4 == 3'h4; // @[RA_Mul.scala 62:44:@436.4]
  assign _T_200 = _T_197 | _T_199; // @[RA_Mul.scala 62:32:@437.4]
  assign _T_203 = io_eB_4 == 3'h1; // @[RA_Mul.scala 64:25:@442.6]
  assign _T_205 = io_eB_4 == 3'h2; // @[RA_Mul.scala 66:25:@447.8]
  assign _T_209 = io_eB_4 == 3'h5; // @[RA_Mul.scala 68:25:@454.10]
  assign _T_212 = io_eB_4 == 3'h6; // @[RA_Mul.scala 70:25:@460.12]
  assign _GEN_20 = _T_212 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@461.12]
  assign _GEN_21 = _T_209 ? _T_106 : _GEN_20; // @[RA_Mul.scala 68:39:@455.10]
  assign _GEN_22 = _T_205 ? _T_103 : _GEN_21; // @[RA_Mul.scala 66:39:@448.8]
  assign _GEN_23 = _T_203 ? io_A : _GEN_22; // @[RA_Mul.scala 64:39:@443.6]
  assign S_v_4 = io_eB_4[2]; // @[RA_Mul.scala 76:23:@470.4]
  assign _T_220 = S_v_4 ^ _T_115; // @[RA_Mul.scala 77:30:@474.4]
  assign SC_v_4 = ~ _T_220; // @[RA_Mul.scala 77:16:@475.4]
  assign _T_223 = io_eB_5 == 3'h0; // @[RA_Mul.scala 62:19:@477.4]
  assign _T_225 = io_eB_5 == 3'h4; // @[RA_Mul.scala 62:44:@478.4]
  assign _T_226 = _T_223 | _T_225; // @[RA_Mul.scala 62:32:@479.4]
  assign _T_229 = io_eB_5 == 3'h1; // @[RA_Mul.scala 64:25:@484.6]
  assign _T_231 = io_eB_5 == 3'h2; // @[RA_Mul.scala 66:25:@489.8]
  assign _T_235 = io_eB_5 == 3'h5; // @[RA_Mul.scala 68:25:@496.10]
  assign _T_238 = io_eB_5 == 3'h6; // @[RA_Mul.scala 70:25:@502.12]
  assign _GEN_25 = _T_238 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@503.12]
  assign _GEN_26 = _T_235 ? _T_106 : _GEN_25; // @[RA_Mul.scala 68:39:@497.10]
  assign _GEN_27 = _T_231 ? _T_103 : _GEN_26; // @[RA_Mul.scala 66:39:@490.8]
  assign _GEN_28 = _T_229 ? io_A : _GEN_27; // @[RA_Mul.scala 64:39:@485.6]
  assign S_v_5 = io_eB_5[2]; // @[RA_Mul.scala 76:23:@512.4]
  assign _T_246 = S_v_5 ^ _T_115; // @[RA_Mul.scala 77:30:@516.4]
  assign SC_v_5 = ~ _T_246; // @[RA_Mul.scala 77:16:@517.4]
  assign _T_249 = io_eB_6 == 3'h0; // @[RA_Mul.scala 62:19:@519.4]
  assign _T_251 = io_eB_6 == 3'h4; // @[RA_Mul.scala 62:44:@520.4]
  assign _T_252 = _T_249 | _T_251; // @[RA_Mul.scala 62:32:@521.4]
  assign _T_255 = io_eB_6 == 3'h1; // @[RA_Mul.scala 64:25:@526.6]
  assign _T_257 = io_eB_6 == 3'h2; // @[RA_Mul.scala 66:25:@531.8]
  assign _T_261 = io_eB_6 == 3'h5; // @[RA_Mul.scala 68:25:@538.10]
  assign _T_264 = io_eB_6 == 3'h6; // @[RA_Mul.scala 70:25:@544.12]
  assign _GEN_30 = _T_264 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@545.12]
  assign _GEN_31 = _T_261 ? _T_106 : _GEN_30; // @[RA_Mul.scala 68:39:@539.10]
  assign _GEN_32 = _T_257 ? _T_103 : _GEN_31; // @[RA_Mul.scala 66:39:@532.8]
  assign _GEN_33 = _T_255 ? io_A : _GEN_32; // @[RA_Mul.scala 64:39:@527.6]
  assign S_v_6 = io_eB_6[2]; // @[RA_Mul.scala 76:23:@554.4]
  assign _T_272 = S_v_6 ^ _T_115; // @[RA_Mul.scala 77:30:@558.4]
  assign SC_v_6 = ~ _T_272; // @[RA_Mul.scala 77:16:@559.4]
  assign _T_275 = io_eB_7 == 3'h0; // @[RA_Mul.scala 62:19:@561.4]
  assign _T_277 = io_eB_7 == 3'h4; // @[RA_Mul.scala 62:44:@562.4]
  assign _T_278 = _T_275 | _T_277; // @[RA_Mul.scala 62:32:@563.4]
  assign _T_281 = io_eB_7 == 3'h1; // @[RA_Mul.scala 64:25:@568.6]
  assign _T_283 = io_eB_7 == 3'h2; // @[RA_Mul.scala 66:25:@573.8]
  assign _T_287 = io_eB_7 == 3'h5; // @[RA_Mul.scala 68:25:@580.10]
  assign _T_290 = io_eB_7 == 3'h6; // @[RA_Mul.scala 70:25:@586.12]
  assign _GEN_35 = _T_290 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@587.12]
  assign _GEN_36 = _T_287 ? _T_106 : _GEN_35; // @[RA_Mul.scala 68:39:@581.10]
  assign _GEN_37 = _T_283 ? _T_103 : _GEN_36; // @[RA_Mul.scala 66:39:@574.8]
  assign _GEN_38 = _T_281 ? io_A : _GEN_37; // @[RA_Mul.scala 64:39:@569.6]
  assign S_v_7 = io_eB_7[2]; // @[RA_Mul.scala 76:23:@596.4]
  assign _T_298 = S_v_7 ^ _T_115; // @[RA_Mul.scala 77:30:@600.4]
  assign SC_v_7 = ~ _T_298; // @[RA_Mul.scala 77:16:@601.4]
  assign _T_300 = {S_v_1,S_v_0}; // @[RA_Mul.scala 79:21:@603.4]
  assign _T_301 = {S_v_3,S_v_2}; // @[RA_Mul.scala 79:21:@604.4]
  assign _T_302 = {_T_301,_T_300}; // @[RA_Mul.scala 79:21:@605.4]
  assign _T_303 = {S_v_5,S_v_4}; // @[RA_Mul.scala 79:21:@606.4]
  assign _T_304 = {S_v_7,S_v_6}; // @[RA_Mul.scala 79:21:@607.4]
  assign _T_305 = {_T_304,_T_303}; // @[RA_Mul.scala 79:21:@608.4]
  assign _T_307 = {SC_v_1,SC_v_0}; // @[RA_Mul.scala 80:23:@611.4]
  assign _T_308 = {SC_v_3,SC_v_2}; // @[RA_Mul.scala 80:23:@612.4]
  assign _T_309 = {_T_308,_T_307}; // @[RA_Mul.scala 80:23:@613.4]
  assign _T_310 = {SC_v_5,SC_v_4}; // @[RA_Mul.scala 80:23:@614.4]
  assign _T_311 = {SC_v_7,SC_v_6}; // @[RA_Mul.scala 80:23:@615.4]
  assign _T_312 = {_T_311,_T_310}; // @[RA_Mul.scala 80:23:@616.4]
  assign io_PP_0 = _T_96 ? 16'h0 : _GEN_3; // @[RA_Mul.scala 63:16:@271.6 RA_Mul.scala 65:16:@276.8 RA_Mul.scala 67:16:@283.10 RA_Mul.scala 69:16:@289.12 RA_Mul.scala 71:16:@297.14 RA_Mul.scala 73:16:@300.14]
  assign io_PP_1 = _T_122 ? 16'h0 : _GEN_8; // @[RA_Mul.scala 63:16:@313.6 RA_Mul.scala 65:16:@318.8 RA_Mul.scala 67:16:@325.10 RA_Mul.scala 69:16:@331.12 RA_Mul.scala 71:16:@339.14 RA_Mul.scala 73:16:@342.14]
  assign io_PP_2 = _T_148 ? 16'h0 : _GEN_13; // @[RA_Mul.scala 63:16:@355.6 RA_Mul.scala 65:16:@360.8 RA_Mul.scala 67:16:@367.10 RA_Mul.scala 69:16:@373.12 RA_Mul.scala 71:16:@381.14 RA_Mul.scala 73:16:@384.14]
  assign io_PP_3 = _T_174 ? 16'h0 : _GEN_18; // @[RA_Mul.scala 63:16:@397.6 RA_Mul.scala 65:16:@402.8 RA_Mul.scala 67:16:@409.10 RA_Mul.scala 69:16:@415.12 RA_Mul.scala 71:16:@423.14 RA_Mul.scala 73:16:@426.14]
  assign io_PP_4 = _T_200 ? 16'h0 : _GEN_23; // @[RA_Mul.scala 63:16:@439.6 RA_Mul.scala 65:16:@444.8 RA_Mul.scala 67:16:@451.10 RA_Mul.scala 69:16:@457.12 RA_Mul.scala 71:16:@465.14 RA_Mul.scala 73:16:@468.14]
  assign io_PP_5 = _T_226 ? 16'h0 : _GEN_28; // @[RA_Mul.scala 63:16:@481.6 RA_Mul.scala 65:16:@486.8 RA_Mul.scala 67:16:@493.10 RA_Mul.scala 69:16:@499.12 RA_Mul.scala 71:16:@507.14 RA_Mul.scala 73:16:@510.14]
  assign io_PP_6 = _T_252 ? 16'h0 : _GEN_33; // @[RA_Mul.scala 63:16:@523.6 RA_Mul.scala 65:16:@528.8 RA_Mul.scala 67:16:@535.10 RA_Mul.scala 69:16:@541.12 RA_Mul.scala 71:16:@549.14 RA_Mul.scala 73:16:@552.14]
  assign io_PP_7 = _T_278 ? 16'h0 : _GEN_38; // @[RA_Mul.scala 63:16:@565.6 RA_Mul.scala 65:16:@570.8 RA_Mul.scala 67:16:@577.10 RA_Mul.scala 69:16:@583.12 RA_Mul.scala 71:16:@591.14 RA_Mul.scala 73:16:@594.14]
  assign io_SC = {_T_312,_T_309}; // @[RA_Mul.scala 80:9:@618.4]
  assign io_S = {_T_305,_T_302}; // @[RA_Mul.scala 79:8:@610.4]
endmodule
module RAMul( // @[:@620.2]
  input         clock, // @[:@621.4]
  input         reset, // @[:@622.4]
  output [15:0] io_PP_0, // @[:@623.4]
  output [15:0] io_PP_1, // @[:@623.4]
  output [15:0] io_PP_2, // @[:@623.4]
  output [15:0] io_PP_3, // @[:@623.4]
  output [15:0] io_PP_4, // @[:@623.4]
  output [15:0] io_PP_5, // @[:@623.4]
  output [15:0] io_PP_6, // @[:@623.4]
  output [15:0] io_PP_7, // @[:@623.4]
  output [15:0] io_SS, // @[:@623.4]
  output [7:0]  io_SC, // @[:@623.4]
  output [7:0]  io_S, // @[:@623.4]
  input  [15:0] io_B, // @[:@623.4]
  input  [15:0] io_A // @[:@623.4]
);
  wire [2:0] BoothEncoder_io_eB_0; // @[RA_Mul.scala 95:28:@625.4]
  wire [2:0] BoothEncoder_io_eB_1; // @[RA_Mul.scala 95:28:@625.4]
  wire [2:0] BoothEncoder_io_eB_2; // @[RA_Mul.scala 95:28:@625.4]
  wire [2:0] BoothEncoder_io_eB_3; // @[RA_Mul.scala 95:28:@625.4]
  wire [2:0] BoothEncoder_io_eB_4; // @[RA_Mul.scala 95:28:@625.4]
  wire [2:0] BoothEncoder_io_eB_5; // @[RA_Mul.scala 95:28:@625.4]
  wire [2:0] BoothEncoder_io_eB_6; // @[RA_Mul.scala 95:28:@625.4]
  wire [2:0] BoothEncoder_io_eB_7; // @[RA_Mul.scala 95:28:@625.4]
  wire [15:0] BoothEncoder_io_B; // @[RA_Mul.scala 95:28:@625.4]
  wire [15:0] PPGenerator_io_PP_0; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_PP_1; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_PP_2; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_PP_3; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_PP_4; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_PP_5; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_PP_6; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_PP_7; // @[RA_Mul.scala 96:27:@628.4]
  wire [7:0] PPGenerator_io_SC; // @[RA_Mul.scala 96:27:@628.4]
  wire [7:0] PPGenerator_io_S; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_0; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_1; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_2; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_3; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_4; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_5; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_6; // @[RA_Mul.scala 96:27:@628.4]
  wire [2:0] PPGenerator_io_eB_7; // @[RA_Mul.scala 96:27:@628.4]
  wire [15:0] PPGenerator_io_A; // @[RA_Mul.scala 96:27:@628.4]
  BoothEncoder_radix4 BoothEncoder ( // @[RA_Mul.scala 95:28:@625.4]
    .io_eB_0(BoothEncoder_io_eB_0),
    .io_eB_1(BoothEncoder_io_eB_1),
    .io_eB_2(BoothEncoder_io_eB_2),
    .io_eB_3(BoothEncoder_io_eB_3),
    .io_eB_4(BoothEncoder_io_eB_4),
    .io_eB_5(BoothEncoder_io_eB_5),
    .io_eB_6(BoothEncoder_io_eB_6),
    .io_eB_7(BoothEncoder_io_eB_7),
    .io_B(BoothEncoder_io_B)
  );
  PPGen PPGenerator ( // @[RA_Mul.scala 96:27:@628.4]
    .io_PP_0(PPGenerator_io_PP_0),
    .io_PP_1(PPGenerator_io_PP_1),
    .io_PP_2(PPGenerator_io_PP_2),
    .io_PP_3(PPGenerator_io_PP_3),
    .io_PP_4(PPGenerator_io_PP_4),
    .io_PP_5(PPGenerator_io_PP_5),
    .io_PP_6(PPGenerator_io_PP_6),
    .io_PP_7(PPGenerator_io_PP_7),
    .io_SC(PPGenerator_io_SC),
    .io_S(PPGenerator_io_S),
    .io_eB_0(PPGenerator_io_eB_0),
    .io_eB_1(PPGenerator_io_eB_1),
    .io_eB_2(PPGenerator_io_eB_2),
    .io_eB_3(PPGenerator_io_eB_3),
    .io_eB_4(PPGenerator_io_eB_4),
    .io_eB_5(PPGenerator_io_eB_5),
    .io_eB_6(PPGenerator_io_eB_6),
    .io_eB_7(PPGenerator_io_eB_7),
    .io_A(PPGenerator_io_A)
  );
  assign io_PP_0 = PPGenerator_io_PP_0; // @[RA_Mul.scala 101:9:@641.4]
  assign io_PP_1 = PPGenerator_io_PP_1; // @[RA_Mul.scala 101:9:@642.4]
  assign io_PP_2 = PPGenerator_io_PP_2; // @[RA_Mul.scala 101:9:@643.4]
  assign io_PP_3 = PPGenerator_io_PP_3; // @[RA_Mul.scala 101:9:@644.4]
  assign io_PP_4 = PPGenerator_io_PP_4; // @[RA_Mul.scala 101:9:@645.4]
  assign io_PP_5 = PPGenerator_io_PP_5; // @[RA_Mul.scala 101:9:@646.4]
  assign io_PP_6 = PPGenerator_io_PP_6; // @[RA_Mul.scala 101:9:@647.4]
  assign io_PP_7 = PPGenerator_io_PP_7; // @[RA_Mul.scala 101:9:@648.4]
  assign io_SS = 16'haaab; // @[RA_Mul.scala 102:9:@649.4]
  assign io_SC = PPGenerator_io_SC; // @[RA_Mul.scala 103:9:@650.4]
  assign io_S = PPGenerator_io_S; // @[RA_Mul.scala 104:8:@651.4]
  assign BoothEncoder_io_B = io_B; // @[RA_Mul.scala 98:21:@631.4]
  assign PPGenerator_io_eB_0 = BoothEncoder_io_eB_0; // @[RA_Mul.scala 99:21:@632.4]
  assign PPGenerator_io_eB_1 = BoothEncoder_io_eB_1; // @[RA_Mul.scala 99:21:@633.4]
  assign PPGenerator_io_eB_2 = BoothEncoder_io_eB_2; // @[RA_Mul.scala 99:21:@634.4]
  assign PPGenerator_io_eB_3 = BoothEncoder_io_eB_3; // @[RA_Mul.scala 99:21:@635.4]
  assign PPGenerator_io_eB_4 = BoothEncoder_io_eB_4; // @[RA_Mul.scala 99:21:@636.4]
  assign PPGenerator_io_eB_5 = BoothEncoder_io_eB_5; // @[RA_Mul.scala 99:21:@637.4]
  assign PPGenerator_io_eB_6 = BoothEncoder_io_eB_6; // @[RA_Mul.scala 99:21:@638.4]
  assign PPGenerator_io_eB_7 = BoothEncoder_io_eB_7; // @[RA_Mul.scala 99:21:@639.4]
  assign PPGenerator_io_A = io_A; // @[RA_Mul.scala 100:20:@640.4]
endmodule
