module HA( // @[:@3.2]
  output  io_s, // @[:@6.4]
  output  io_cout, // @[:@6.4]
  input   io_a, // @[:@6.4]
  input   io_b // @[:@6.4]
);
  assign io_s = io_a ^ io_b; // @[RA_Mul.scala 12:8:@11.4]
  assign io_cout = io_a & io_b; // @[RA_Mul.scala 11:11:@9.4]
endmodule
module FA( // @[:@13.2]
  output  io_s, // @[:@16.4]
  output  io_cout, // @[:@16.4]
  input   io_a, // @[:@16.4]
  input   io_b, // @[:@16.4]
  input   io_cin // @[:@16.4]
);
  wire  _T_15; // @[RA_Mul.scala 35:16:@18.4]
  wire  _T_17; // @[RA_Mul.scala 36:20:@21.4]
  wire  _T_18; // @[RA_Mul.scala 36:36:@22.4]
  wire  _T_19; // @[RA_Mul.scala 36:28:@23.4]
  wire  _T_20; // @[RA_Mul.scala 36:54:@24.4]
  assign _T_15 = io_a ^ io_b; // @[RA_Mul.scala 35:16:@18.4]
  assign _T_17 = io_a & io_b; // @[RA_Mul.scala 36:20:@21.4]
  assign _T_18 = io_a & io_cin; // @[RA_Mul.scala 36:36:@22.4]
  assign _T_19 = _T_17 | _T_18; // @[RA_Mul.scala 36:28:@23.4]
  assign _T_20 = io_b & io_cin; // @[RA_Mul.scala 36:54:@24.4]
  assign io_s = _T_15 ^ io_cin; // @[RA_Mul.scala 35:8:@20.4]
  assign io_cout = _T_19 | _T_20; // @[RA_Mul.scala 36:11:@26.4]
endmodule
module Reduction_3( // @[:@298.2]
  input   clock, // @[:@299.4]
  input   reset, // @[:@300.4]
  output  io_matrix_o_0_0, // @[:@301.4]
  output  io_matrix_o_0_1, // @[:@301.4]
  output  io_matrix_o_0_2, // @[:@301.4]
  output  io_matrix_o_0_3, // @[:@301.4]
  output  io_matrix_o_0_4, // @[:@301.4]
  output  io_matrix_o_0_5, // @[:@301.4]
  output  io_matrix_o_0_6, // @[:@301.4]
  output  io_matrix_o_0_7, // @[:@301.4]
  output  io_matrix_o_0_8, // @[:@301.4]
  output  io_matrix_o_0_9, // @[:@301.4]
  output  io_matrix_o_0_10, // @[:@301.4]
  output  io_matrix_o_0_11, // @[:@301.4]
  output  io_matrix_o_0_12, // @[:@301.4]
  output  io_matrix_o_0_13, // @[:@301.4]
  output  io_matrix_o_0_14, // @[:@301.4]
  output  io_matrix_o_0_15, // @[:@301.4]
  output  io_matrix_o_0_16, // @[:@301.4]
  output  io_matrix_o_0_17, // @[:@301.4]
  output  io_matrix_o_0_18, // @[:@301.4]
  output  io_matrix_o_0_19, // @[:@301.4]
  output  io_matrix_o_0_20, // @[:@301.4]
  output  io_matrix_o_0_21, // @[:@301.4]
  output  io_matrix_o_0_22, // @[:@301.4]
  output  io_matrix_o_0_23, // @[:@301.4]
  output  io_matrix_o_0_24, // @[:@301.4]
  output  io_matrix_o_0_25, // @[:@301.4]
  output  io_matrix_o_0_26, // @[:@301.4]
  output  io_matrix_o_0_27, // @[:@301.4]
  output  io_matrix_o_0_28, // @[:@301.4]
  output  io_matrix_o_0_29, // @[:@301.4]
  output  io_matrix_o_0_30, // @[:@301.4]
  output  io_matrix_o_0_31, // @[:@301.4]
  output  io_matrix_o_1_0, // @[:@301.4]
  output  io_matrix_o_1_1, // @[:@301.4]
  output  io_matrix_o_1_2, // @[:@301.4]
  output  io_matrix_o_1_3, // @[:@301.4]
  output  io_matrix_o_1_4, // @[:@301.4]
  output  io_matrix_o_1_5, // @[:@301.4]
  output  io_matrix_o_1_6, // @[:@301.4]
  output  io_matrix_o_1_7, // @[:@301.4]
  output  io_matrix_o_1_8, // @[:@301.4]
  output  io_matrix_o_1_9, // @[:@301.4]
  output  io_matrix_o_1_10, // @[:@301.4]
  output  io_matrix_o_1_11, // @[:@301.4]
  output  io_matrix_o_1_12, // @[:@301.4]
  output  io_matrix_o_1_13, // @[:@301.4]
  output  io_matrix_o_1_14, // @[:@301.4]
  output  io_matrix_o_1_15, // @[:@301.4]
  output  io_matrix_o_1_16, // @[:@301.4]
  output  io_matrix_o_1_17, // @[:@301.4]
  output  io_matrix_o_1_18, // @[:@301.4]
  output  io_matrix_o_1_19, // @[:@301.4]
  output  io_matrix_o_1_20, // @[:@301.4]
  output  io_matrix_o_1_21, // @[:@301.4]
  output  io_matrix_o_1_22, // @[:@301.4]
  output  io_matrix_o_1_23, // @[:@301.4]
  output  io_matrix_o_1_24, // @[:@301.4]
  output  io_matrix_o_1_25, // @[:@301.4]
  output  io_matrix_o_1_26, // @[:@301.4]
  output  io_matrix_o_1_27, // @[:@301.4]
  output  io_matrix_o_1_28, // @[:@301.4]
  output  io_matrix_o_1_29, // @[:@301.4]
  output  io_matrix_o_1_30, // @[:@301.4]
  output  io_matrix_o_1_31, // @[:@301.4]
  output  io_matrix_o_2_0, // @[:@301.4]
  output  io_matrix_o_2_1, // @[:@301.4]
  output  io_matrix_o_2_2, // @[:@301.4]
  output  io_matrix_o_2_3, // @[:@301.4]
  output  io_matrix_o_2_4, // @[:@301.4]
  output  io_matrix_o_2_5, // @[:@301.4]
  output  io_matrix_o_2_6, // @[:@301.4]
  output  io_matrix_o_2_7, // @[:@301.4]
  output  io_matrix_o_2_8, // @[:@301.4]
  output  io_matrix_o_2_9, // @[:@301.4]
  output  io_matrix_o_2_10, // @[:@301.4]
  output  io_matrix_o_2_11, // @[:@301.4]
  output  io_matrix_o_2_12, // @[:@301.4]
  output  io_matrix_o_2_13, // @[:@301.4]
  output  io_matrix_o_2_14, // @[:@301.4]
  output  io_matrix_o_2_15, // @[:@301.4]
  output  io_matrix_o_2_16, // @[:@301.4]
  output  io_matrix_o_2_17, // @[:@301.4]
  output  io_matrix_o_2_18, // @[:@301.4]
  output  io_matrix_o_2_19, // @[:@301.4]
  output  io_matrix_o_2_20, // @[:@301.4]
  output  io_matrix_o_2_21, // @[:@301.4]
  output  io_matrix_o_2_22, // @[:@301.4]
  output  io_matrix_o_2_23, // @[:@301.4]
  output  io_matrix_o_2_24, // @[:@301.4]
  output  io_matrix_o_2_25, // @[:@301.4]
  output  io_matrix_o_2_26, // @[:@301.4]
  output  io_matrix_o_2_27, // @[:@301.4]
  output  io_matrix_o_2_28, // @[:@301.4]
  output  io_matrix_o_2_29, // @[:@301.4]
  output  io_matrix_o_2_30, // @[:@301.4]
  output  io_matrix_o_2_31, // @[:@301.4]
  input   io_matrix_i_0_0, // @[:@301.4]
  input   io_matrix_i_0_1, // @[:@301.4]
  input   io_matrix_i_0_2, // @[:@301.4]
  input   io_matrix_i_0_3, // @[:@301.4]
  input   io_matrix_i_0_4, // @[:@301.4]
  input   io_matrix_i_0_5, // @[:@301.4]
  input   io_matrix_i_0_6, // @[:@301.4]
  input   io_matrix_i_0_7, // @[:@301.4]
  input   io_matrix_i_0_8, // @[:@301.4]
  input   io_matrix_i_0_9, // @[:@301.4]
  input   io_matrix_i_0_10, // @[:@301.4]
  input   io_matrix_i_0_11, // @[:@301.4]
  input   io_matrix_i_0_12, // @[:@301.4]
  input   io_matrix_i_0_13, // @[:@301.4]
  input   io_matrix_i_0_14, // @[:@301.4]
  input   io_matrix_i_0_15, // @[:@301.4]
  input   io_matrix_i_0_16, // @[:@301.4]
  input   io_matrix_i_0_17, // @[:@301.4]
  input   io_matrix_i_0_18, // @[:@301.4]
  input   io_matrix_i_0_19, // @[:@301.4]
  input   io_matrix_i_0_20, // @[:@301.4]
  input   io_matrix_i_0_21, // @[:@301.4]
  input   io_matrix_i_0_22, // @[:@301.4]
  input   io_matrix_i_0_23, // @[:@301.4]
  input   io_matrix_i_0_24, // @[:@301.4]
  input   io_matrix_i_0_25, // @[:@301.4]
  input   io_matrix_i_0_26, // @[:@301.4]
  input   io_matrix_i_0_27, // @[:@301.4]
  input   io_matrix_i_0_28, // @[:@301.4]
  input   io_matrix_i_0_29, // @[:@301.4]
  input   io_matrix_i_0_30, // @[:@301.4]
  input   io_matrix_i_0_31, // @[:@301.4]
  input   io_matrix_i_1_0, // @[:@301.4]
  input   io_matrix_i_1_1, // @[:@301.4]
  input   io_matrix_i_1_2, // @[:@301.4]
  input   io_matrix_i_1_3, // @[:@301.4]
  input   io_matrix_i_1_4, // @[:@301.4]
  input   io_matrix_i_1_5, // @[:@301.4]
  input   io_matrix_i_1_6, // @[:@301.4]
  input   io_matrix_i_1_7, // @[:@301.4]
  input   io_matrix_i_1_8, // @[:@301.4]
  input   io_matrix_i_1_9, // @[:@301.4]
  input   io_matrix_i_1_10, // @[:@301.4]
  input   io_matrix_i_1_11, // @[:@301.4]
  input   io_matrix_i_1_12, // @[:@301.4]
  input   io_matrix_i_1_13, // @[:@301.4]
  input   io_matrix_i_1_14, // @[:@301.4]
  input   io_matrix_i_1_15, // @[:@301.4]
  input   io_matrix_i_1_16, // @[:@301.4]
  input   io_matrix_i_1_17, // @[:@301.4]
  input   io_matrix_i_1_18, // @[:@301.4]
  input   io_matrix_i_1_19, // @[:@301.4]
  input   io_matrix_i_1_20, // @[:@301.4]
  input   io_matrix_i_1_21, // @[:@301.4]
  input   io_matrix_i_1_22, // @[:@301.4]
  input   io_matrix_i_1_23, // @[:@301.4]
  input   io_matrix_i_1_24, // @[:@301.4]
  input   io_matrix_i_1_25, // @[:@301.4]
  input   io_matrix_i_1_26, // @[:@301.4]
  input   io_matrix_i_1_27, // @[:@301.4]
  input   io_matrix_i_1_28, // @[:@301.4]
  input   io_matrix_i_1_29, // @[:@301.4]
  input   io_matrix_i_1_30, // @[:@301.4]
  input   io_matrix_i_1_31, // @[:@301.4]
  input   io_matrix_i_2_0, // @[:@301.4]
  input   io_matrix_i_2_1, // @[:@301.4]
  input   io_matrix_i_2_2, // @[:@301.4]
  input   io_matrix_i_2_3, // @[:@301.4]
  input   io_matrix_i_2_4, // @[:@301.4]
  input   io_matrix_i_2_5, // @[:@301.4]
  input   io_matrix_i_2_6, // @[:@301.4]
  input   io_matrix_i_2_7, // @[:@301.4]
  input   io_matrix_i_2_8, // @[:@301.4]
  input   io_matrix_i_2_9, // @[:@301.4]
  input   io_matrix_i_2_10, // @[:@301.4]
  input   io_matrix_i_2_11, // @[:@301.4]
  input   io_matrix_i_2_12, // @[:@301.4]
  input   io_matrix_i_2_13, // @[:@301.4]
  input   io_matrix_i_2_14, // @[:@301.4]
  input   io_matrix_i_2_15, // @[:@301.4]
  input   io_matrix_i_2_16, // @[:@301.4]
  input   io_matrix_i_2_17, // @[:@301.4]
  input   io_matrix_i_2_18, // @[:@301.4]
  input   io_matrix_i_2_19, // @[:@301.4]
  input   io_matrix_i_2_20, // @[:@301.4]
  input   io_matrix_i_2_21, // @[:@301.4]
  input   io_matrix_i_2_22, // @[:@301.4]
  input   io_matrix_i_2_23, // @[:@301.4]
  input   io_matrix_i_2_24, // @[:@301.4]
  input   io_matrix_i_2_25, // @[:@301.4]
  input   io_matrix_i_2_26, // @[:@301.4]
  input   io_matrix_i_2_27, // @[:@301.4]
  input   io_matrix_i_2_28, // @[:@301.4]
  input   io_matrix_i_2_29, // @[:@301.4]
  input   io_matrix_i_2_30, // @[:@301.4]
  input   io_matrix_i_2_31, // @[:@301.4]
  input   io_matrix_i_3_0, // @[:@301.4]
  input   io_matrix_i_3_1, // @[:@301.4]
  input   io_matrix_i_3_2, // @[:@301.4]
  input   io_matrix_i_3_3, // @[:@301.4]
  input   io_matrix_i_3_4, // @[:@301.4]
  input   io_matrix_i_3_5, // @[:@301.4]
  input   io_matrix_i_3_6, // @[:@301.4]
  input   io_matrix_i_3_7, // @[:@301.4]
  input   io_matrix_i_3_8, // @[:@301.4]
  input   io_matrix_i_3_9, // @[:@301.4]
  input   io_matrix_i_3_10, // @[:@301.4]
  input   io_matrix_i_3_11, // @[:@301.4]
  input   io_matrix_i_3_12, // @[:@301.4]
  input   io_matrix_i_3_13, // @[:@301.4]
  input   io_matrix_i_3_14, // @[:@301.4]
  input   io_matrix_i_3_15, // @[:@301.4]
  input   io_matrix_i_3_16, // @[:@301.4]
  input   io_matrix_i_3_17, // @[:@301.4]
  input   io_matrix_i_3_18, // @[:@301.4]
  input   io_matrix_i_3_19, // @[:@301.4]
  input   io_matrix_i_3_20, // @[:@301.4]
  input   io_matrix_i_3_21, // @[:@301.4]
  input   io_matrix_i_3_22, // @[:@301.4]
  input   io_matrix_i_3_23, // @[:@301.4]
  input   io_matrix_i_3_24, // @[:@301.4]
  input   io_matrix_i_3_25, // @[:@301.4]
  input   io_matrix_i_3_26, // @[:@301.4]
  input   io_matrix_i_3_27, // @[:@301.4]
  input   io_matrix_i_3_28, // @[:@301.4]
  input   io_matrix_i_3_29, // @[:@301.4]
  input   io_matrix_i_3_30, // @[:@301.4]
  input   io_matrix_i_3_31 // @[:@301.4]
);
  wire  HA_io_s; // @[RA_Mul.scala 18:21:@309.4]
  wire  HA_io_cout; // @[RA_Mul.scala 18:21:@309.4]
  wire  HA_io_a; // @[RA_Mul.scala 18:21:@309.4]
  wire  HA_io_b; // @[RA_Mul.scala 18:21:@309.4]
  wire  FA_io_s; // @[RA_Mul.scala 42:21:@320.4]
  wire  FA_io_cout; // @[RA_Mul.scala 42:21:@320.4]
  wire  FA_io_a; // @[RA_Mul.scala 42:21:@320.4]
  wire  FA_io_b; // @[RA_Mul.scala 42:21:@320.4]
  wire  FA_io_cin; // @[RA_Mul.scala 42:21:@320.4]
  wire  FA_1_io_s; // @[RA_Mul.scala 42:21:@341.4]
  wire  FA_1_io_cout; // @[RA_Mul.scala 42:21:@341.4]
  wire  FA_1_io_a; // @[RA_Mul.scala 42:21:@341.4]
  wire  FA_1_io_b; // @[RA_Mul.scala 42:21:@341.4]
  wire  FA_1_io_cin; // @[RA_Mul.scala 42:21:@341.4]
  wire  FA_2_io_s; // @[RA_Mul.scala 42:21:@351.4]
  wire  FA_2_io_cout; // @[RA_Mul.scala 42:21:@351.4]
  wire  FA_2_io_a; // @[RA_Mul.scala 42:21:@351.4]
  wire  FA_2_io_b; // @[RA_Mul.scala 42:21:@351.4]
  wire  FA_2_io_cin; // @[RA_Mul.scala 42:21:@351.4]
  wire  FA_3_io_s; // @[RA_Mul.scala 42:21:@360.4]
  wire  FA_3_io_cout; // @[RA_Mul.scala 42:21:@360.4]
  wire  FA_3_io_a; // @[RA_Mul.scala 42:21:@360.4]
  wire  FA_3_io_b; // @[RA_Mul.scala 42:21:@360.4]
  wire  FA_3_io_cin; // @[RA_Mul.scala 42:21:@360.4]
  wire  FA_4_io_s; // @[RA_Mul.scala 42:21:@369.4]
  wire  FA_4_io_cout; // @[RA_Mul.scala 42:21:@369.4]
  wire  FA_4_io_a; // @[RA_Mul.scala 42:21:@369.4]
  wire  FA_4_io_b; // @[RA_Mul.scala 42:21:@369.4]
  wire  FA_4_io_cin; // @[RA_Mul.scala 42:21:@369.4]
  wire  FA_5_io_s; // @[RA_Mul.scala 42:21:@378.4]
  wire  FA_5_io_cout; // @[RA_Mul.scala 42:21:@378.4]
  wire  FA_5_io_a; // @[RA_Mul.scala 42:21:@378.4]
  wire  FA_5_io_b; // @[RA_Mul.scala 42:21:@378.4]
  wire  FA_5_io_cin; // @[RA_Mul.scala 42:21:@378.4]
  wire  FA_6_io_s; // @[RA_Mul.scala 42:21:@387.4]
  wire  FA_6_io_cout; // @[RA_Mul.scala 42:21:@387.4]
  wire  FA_6_io_a; // @[RA_Mul.scala 42:21:@387.4]
  wire  FA_6_io_b; // @[RA_Mul.scala 42:21:@387.4]
  wire  FA_6_io_cin; // @[RA_Mul.scala 42:21:@387.4]
  wire  FA_7_io_s; // @[RA_Mul.scala 42:21:@396.4]
  wire  FA_7_io_cout; // @[RA_Mul.scala 42:21:@396.4]
  wire  FA_7_io_a; // @[RA_Mul.scala 42:21:@396.4]
  wire  FA_7_io_b; // @[RA_Mul.scala 42:21:@396.4]
  wire  FA_7_io_cin; // @[RA_Mul.scala 42:21:@396.4]
  wire  FA_8_io_s; // @[RA_Mul.scala 42:21:@405.4]
  wire  FA_8_io_cout; // @[RA_Mul.scala 42:21:@405.4]
  wire  FA_8_io_a; // @[RA_Mul.scala 42:21:@405.4]
  wire  FA_8_io_b; // @[RA_Mul.scala 42:21:@405.4]
  wire  FA_8_io_cin; // @[RA_Mul.scala 42:21:@405.4]
  wire  FA_9_io_s; // @[RA_Mul.scala 42:21:@414.4]
  wire  FA_9_io_cout; // @[RA_Mul.scala 42:21:@414.4]
  wire  FA_9_io_a; // @[RA_Mul.scala 42:21:@414.4]
  wire  FA_9_io_b; // @[RA_Mul.scala 42:21:@414.4]
  wire  FA_9_io_cin; // @[RA_Mul.scala 42:21:@414.4]
  wire  FA_10_io_s; // @[RA_Mul.scala 42:21:@423.4]
  wire  FA_10_io_cout; // @[RA_Mul.scala 42:21:@423.4]
  wire  FA_10_io_a; // @[RA_Mul.scala 42:21:@423.4]
  wire  FA_10_io_b; // @[RA_Mul.scala 42:21:@423.4]
  wire  FA_10_io_cin; // @[RA_Mul.scala 42:21:@423.4]
  wire  FA_11_io_s; // @[RA_Mul.scala 42:21:@432.4]
  wire  FA_11_io_cout; // @[RA_Mul.scala 42:21:@432.4]
  wire  FA_11_io_a; // @[RA_Mul.scala 42:21:@432.4]
  wire  FA_11_io_b; // @[RA_Mul.scala 42:21:@432.4]
  wire  FA_11_io_cin; // @[RA_Mul.scala 42:21:@432.4]
  wire  FA_12_io_s; // @[RA_Mul.scala 42:21:@441.4]
  wire  FA_12_io_cout; // @[RA_Mul.scala 42:21:@441.4]
  wire  FA_12_io_a; // @[RA_Mul.scala 42:21:@441.4]
  wire  FA_12_io_b; // @[RA_Mul.scala 42:21:@441.4]
  wire  FA_12_io_cin; // @[RA_Mul.scala 42:21:@441.4]
  wire  FA_13_io_s; // @[RA_Mul.scala 42:21:@450.4]
  wire  FA_13_io_cout; // @[RA_Mul.scala 42:21:@450.4]
  wire  FA_13_io_a; // @[RA_Mul.scala 42:21:@450.4]
  wire  FA_13_io_b; // @[RA_Mul.scala 42:21:@450.4]
  wire  FA_13_io_cin; // @[RA_Mul.scala 42:21:@450.4]
  wire  FA_14_io_s; // @[RA_Mul.scala 42:21:@459.4]
  wire  FA_14_io_cout; // @[RA_Mul.scala 42:21:@459.4]
  wire  FA_14_io_a; // @[RA_Mul.scala 42:21:@459.4]
  wire  FA_14_io_b; // @[RA_Mul.scala 42:21:@459.4]
  wire  FA_14_io_cin; // @[RA_Mul.scala 42:21:@459.4]
  wire  FA_15_io_s; // @[RA_Mul.scala 42:21:@468.4]
  wire  FA_15_io_cout; // @[RA_Mul.scala 42:21:@468.4]
  wire  FA_15_io_a; // @[RA_Mul.scala 42:21:@468.4]
  wire  FA_15_io_b; // @[RA_Mul.scala 42:21:@468.4]
  wire  FA_15_io_cin; // @[RA_Mul.scala 42:21:@468.4]
  wire  FA_16_io_s; // @[RA_Mul.scala 42:21:@477.4]
  wire  FA_16_io_cout; // @[RA_Mul.scala 42:21:@477.4]
  wire  FA_16_io_a; // @[RA_Mul.scala 42:21:@477.4]
  wire  FA_16_io_b; // @[RA_Mul.scala 42:21:@477.4]
  wire  FA_16_io_cin; // @[RA_Mul.scala 42:21:@477.4]
  wire  FA_17_io_s; // @[RA_Mul.scala 42:21:@491.4]
  wire  FA_17_io_cout; // @[RA_Mul.scala 42:21:@491.4]
  wire  FA_17_io_a; // @[RA_Mul.scala 42:21:@491.4]
  wire  FA_17_io_b; // @[RA_Mul.scala 42:21:@491.4]
  wire  FA_17_io_cin; // @[RA_Mul.scala 42:21:@491.4]
  wire  FA_18_io_s; // @[RA_Mul.scala 42:21:@506.4]
  wire  FA_18_io_cout; // @[RA_Mul.scala 42:21:@506.4]
  wire  FA_18_io_a; // @[RA_Mul.scala 42:21:@506.4]
  wire  FA_18_io_b; // @[RA_Mul.scala 42:21:@506.4]
  wire  FA_18_io_cin; // @[RA_Mul.scala 42:21:@506.4]
  HA HA ( // @[RA_Mul.scala 18:21:@309.4]
    .io_s(HA_io_s),
    .io_cout(HA_io_cout),
    .io_a(HA_io_a),
    .io_b(HA_io_b)
  );
  FA FA ( // @[RA_Mul.scala 42:21:@320.4]
    .io_s(FA_io_s),
    .io_cout(FA_io_cout),
    .io_a(FA_io_a),
    .io_b(FA_io_b),
    .io_cin(FA_io_cin)
  );
  FA FA_1 ( // @[RA_Mul.scala 42:21:@341.4]
    .io_s(FA_1_io_s),
    .io_cout(FA_1_io_cout),
    .io_a(FA_1_io_a),
    .io_b(FA_1_io_b),
    .io_cin(FA_1_io_cin)
  );
  FA FA_2 ( // @[RA_Mul.scala 42:21:@351.4]
    .io_s(FA_2_io_s),
    .io_cout(FA_2_io_cout),
    .io_a(FA_2_io_a),
    .io_b(FA_2_io_b),
    .io_cin(FA_2_io_cin)
  );
  FA FA_3 ( // @[RA_Mul.scala 42:21:@360.4]
    .io_s(FA_3_io_s),
    .io_cout(FA_3_io_cout),
    .io_a(FA_3_io_a),
    .io_b(FA_3_io_b),
    .io_cin(FA_3_io_cin)
  );
  FA FA_4 ( // @[RA_Mul.scala 42:21:@369.4]
    .io_s(FA_4_io_s),
    .io_cout(FA_4_io_cout),
    .io_a(FA_4_io_a),
    .io_b(FA_4_io_b),
    .io_cin(FA_4_io_cin)
  );
  FA FA_5 ( // @[RA_Mul.scala 42:21:@378.4]
    .io_s(FA_5_io_s),
    .io_cout(FA_5_io_cout),
    .io_a(FA_5_io_a),
    .io_b(FA_5_io_b),
    .io_cin(FA_5_io_cin)
  );
  FA FA_6 ( // @[RA_Mul.scala 42:21:@387.4]
    .io_s(FA_6_io_s),
    .io_cout(FA_6_io_cout),
    .io_a(FA_6_io_a),
    .io_b(FA_6_io_b),
    .io_cin(FA_6_io_cin)
  );
  FA FA_7 ( // @[RA_Mul.scala 42:21:@396.4]
    .io_s(FA_7_io_s),
    .io_cout(FA_7_io_cout),
    .io_a(FA_7_io_a),
    .io_b(FA_7_io_b),
    .io_cin(FA_7_io_cin)
  );
  FA FA_8 ( // @[RA_Mul.scala 42:21:@405.4]
    .io_s(FA_8_io_s),
    .io_cout(FA_8_io_cout),
    .io_a(FA_8_io_a),
    .io_b(FA_8_io_b),
    .io_cin(FA_8_io_cin)
  );
  FA FA_9 ( // @[RA_Mul.scala 42:21:@414.4]
    .io_s(FA_9_io_s),
    .io_cout(FA_9_io_cout),
    .io_a(FA_9_io_a),
    .io_b(FA_9_io_b),
    .io_cin(FA_9_io_cin)
  );
  FA FA_10 ( // @[RA_Mul.scala 42:21:@423.4]
    .io_s(FA_10_io_s),
    .io_cout(FA_10_io_cout),
    .io_a(FA_10_io_a),
    .io_b(FA_10_io_b),
    .io_cin(FA_10_io_cin)
  );
  FA FA_11 ( // @[RA_Mul.scala 42:21:@432.4]
    .io_s(FA_11_io_s),
    .io_cout(FA_11_io_cout),
    .io_a(FA_11_io_a),
    .io_b(FA_11_io_b),
    .io_cin(FA_11_io_cin)
  );
  FA FA_12 ( // @[RA_Mul.scala 42:21:@441.4]
    .io_s(FA_12_io_s),
    .io_cout(FA_12_io_cout),
    .io_a(FA_12_io_a),
    .io_b(FA_12_io_b),
    .io_cin(FA_12_io_cin)
  );
  FA FA_13 ( // @[RA_Mul.scala 42:21:@450.4]
    .io_s(FA_13_io_s),
    .io_cout(FA_13_io_cout),
    .io_a(FA_13_io_a),
    .io_b(FA_13_io_b),
    .io_cin(FA_13_io_cin)
  );
  FA FA_14 ( // @[RA_Mul.scala 42:21:@459.4]
    .io_s(FA_14_io_s),
    .io_cout(FA_14_io_cout),
    .io_a(FA_14_io_a),
    .io_b(FA_14_io_b),
    .io_cin(FA_14_io_cin)
  );
  FA FA_15 ( // @[RA_Mul.scala 42:21:@468.4]
    .io_s(FA_15_io_s),
    .io_cout(FA_15_io_cout),
    .io_a(FA_15_io_a),
    .io_b(FA_15_io_b),
    .io_cin(FA_15_io_cin)
  );
  FA FA_16 ( // @[RA_Mul.scala 42:21:@477.4]
    .io_s(FA_16_io_s),
    .io_cout(FA_16_io_cout),
    .io_a(FA_16_io_a),
    .io_b(FA_16_io_b),
    .io_cin(FA_16_io_cin)
  );
  FA FA_17 ( // @[RA_Mul.scala 42:21:@491.4]
    .io_s(FA_17_io_s),
    .io_cout(FA_17_io_cout),
    .io_a(FA_17_io_a),
    .io_b(FA_17_io_b),
    .io_cin(FA_17_io_cin)
  );
  FA FA_18 ( // @[RA_Mul.scala 42:21:@506.4]
    .io_s(FA_18_io_s),
    .io_cout(FA_18_io_cout),
    .io_a(FA_18_io_a),
    .io_b(FA_18_io_b),
    .io_cin(FA_18_io_cin)
  );
  assign io_matrix_o_0_0 = io_matrix_i_0_0; // @[RA_Mul.scala 421:21:@303.4]
  assign io_matrix_o_0_1 = io_matrix_i_0_1; // @[RA_Mul.scala 424:21:@306.4]
  assign io_matrix_o_0_2 = HA_io_s; // @[RA_Mul.scala 21:7:@314.4]
  assign io_matrix_o_0_3 = io_matrix_i_0_3; // @[RA_Mul.scala 430:21:@318.4]
  assign io_matrix_o_0_4 = FA_io_s; // @[RA_Mul.scala 46:7:@326.4]
  assign io_matrix_o_0_5 = io_matrix_i_0_5; // @[RA_Mul.scala 436:21:@330.4]
  assign io_matrix_o_0_6 = io_matrix_i_0_6; // @[RA_Mul.scala 440:23:@332.4]
  assign io_matrix_o_0_7 = io_matrix_i_0_7; // @[RA_Mul.scala 440:23:@335.4]
  assign io_matrix_o_0_8 = io_matrix_i_0_8; // @[RA_Mul.scala 440:23:@338.4]
  assign io_matrix_o_0_9 = FA_1_io_s; // @[RA_Mul.scala 46:7:@347.4]
  assign io_matrix_o_0_10 = FA_2_io_s; // @[RA_Mul.scala 46:7:@357.4]
  assign io_matrix_o_0_11 = FA_3_io_s; // @[RA_Mul.scala 46:7:@366.4]
  assign io_matrix_o_0_12 = FA_4_io_s; // @[RA_Mul.scala 46:7:@375.4]
  assign io_matrix_o_0_13 = FA_5_io_s; // @[RA_Mul.scala 46:7:@384.4]
  assign io_matrix_o_0_14 = FA_6_io_s; // @[RA_Mul.scala 46:7:@393.4]
  assign io_matrix_o_0_15 = FA_7_io_s; // @[RA_Mul.scala 46:7:@402.4]
  assign io_matrix_o_0_16 = FA_8_io_s; // @[RA_Mul.scala 46:7:@411.4]
  assign io_matrix_o_0_17 = FA_9_io_s; // @[RA_Mul.scala 46:7:@420.4]
  assign io_matrix_o_0_18 = FA_10_io_s; // @[RA_Mul.scala 46:7:@429.4]
  assign io_matrix_o_0_19 = FA_11_io_s; // @[RA_Mul.scala 46:7:@438.4]
  assign io_matrix_o_0_20 = FA_12_io_s; // @[RA_Mul.scala 46:7:@447.4]
  assign io_matrix_o_0_21 = FA_13_io_s; // @[RA_Mul.scala 46:7:@456.4]
  assign io_matrix_o_0_22 = FA_14_io_s; // @[RA_Mul.scala 46:7:@465.4]
  assign io_matrix_o_0_23 = FA_15_io_s; // @[RA_Mul.scala 46:7:@474.4]
  assign io_matrix_o_0_24 = FA_16_io_s; // @[RA_Mul.scala 46:7:@483.4]
  assign io_matrix_o_0_25 = io_matrix_i_0_25; // @[RA_Mul.scala 468:22:@486.4]
  assign io_matrix_o_0_26 = io_matrix_i_0_26; // @[RA_Mul.scala 471:22:@488.4]
  assign io_matrix_o_0_27 = FA_17_io_s; // @[RA_Mul.scala 46:7:@497.4]
  assign io_matrix_o_0_28 = io_matrix_i_0_28; // @[RA_Mul.scala 478:22:@501.4]
  assign io_matrix_o_0_29 = io_matrix_i_0_29; // @[RA_Mul.scala 481:22:@503.4]
  assign io_matrix_o_0_30 = FA_18_io_s; // @[RA_Mul.scala 46:7:@512.4]
  assign io_matrix_o_0_31 = io_matrix_i_0_31; // @[RA_Mul.scala 487:22:@516.4]
  assign io_matrix_o_1_0 = 1'h0; // @[RA_Mul.scala 417:19:@304.4]
  assign io_matrix_o_1_1 = 1'h0; // @[RA_Mul.scala 417:19:@307.4]
  assign io_matrix_o_1_2 = 1'h0; // @[RA_Mul.scala 417:19:@316.4]
  assign io_matrix_o_1_3 = HA_io_cout; // @[RA_Mul.scala 22:10:@315.4]
  assign io_matrix_o_1_4 = 1'h0; // @[RA_Mul.scala 417:19:@328.4]
  assign io_matrix_o_1_5 = FA_io_cout; // @[RA_Mul.scala 47:10:@327.4]
  assign io_matrix_o_1_6 = io_matrix_i_1_6; // @[RA_Mul.scala 441:23:@333.4]
  assign io_matrix_o_1_7 = io_matrix_i_1_7; // @[RA_Mul.scala 441:23:@336.4]
  assign io_matrix_o_1_8 = io_matrix_i_1_8; // @[RA_Mul.scala 441:23:@339.4]
  assign io_matrix_o_1_9 = io_matrix_i_3_9; // @[RA_Mul.scala 446:21:@349.4]
  assign io_matrix_o_1_10 = FA_1_io_cout; // @[RA_Mul.scala 47:10:@348.4]
  assign io_matrix_o_1_11 = FA_2_io_cout; // @[RA_Mul.scala 47:10:@358.4]
  assign io_matrix_o_1_12 = FA_3_io_cout; // @[RA_Mul.scala 47:10:@367.4]
  assign io_matrix_o_1_13 = FA_4_io_cout; // @[RA_Mul.scala 47:10:@376.4]
  assign io_matrix_o_1_14 = FA_5_io_cout; // @[RA_Mul.scala 47:10:@385.4]
  assign io_matrix_o_1_15 = FA_6_io_cout; // @[RA_Mul.scala 47:10:@394.4]
  assign io_matrix_o_1_16 = FA_7_io_cout; // @[RA_Mul.scala 47:10:@403.4]
  assign io_matrix_o_1_17 = FA_8_io_cout; // @[RA_Mul.scala 47:10:@412.4]
  assign io_matrix_o_1_18 = FA_9_io_cout; // @[RA_Mul.scala 47:10:@421.4]
  assign io_matrix_o_1_19 = FA_10_io_cout; // @[RA_Mul.scala 47:10:@430.4]
  assign io_matrix_o_1_20 = FA_11_io_cout; // @[RA_Mul.scala 47:10:@439.4]
  assign io_matrix_o_1_21 = FA_12_io_cout; // @[RA_Mul.scala 47:10:@448.4]
  assign io_matrix_o_1_22 = FA_13_io_cout; // @[RA_Mul.scala 47:10:@457.4]
  assign io_matrix_o_1_23 = FA_14_io_cout; // @[RA_Mul.scala 47:10:@466.4]
  assign io_matrix_o_1_24 = FA_15_io_cout; // @[RA_Mul.scala 47:10:@475.4]
  assign io_matrix_o_1_25 = FA_16_io_cout; // @[RA_Mul.scala 47:10:@484.4]
  assign io_matrix_o_1_26 = io_matrix_i_1_26; // @[RA_Mul.scala 472:22:@489.4]
  assign io_matrix_o_1_27 = 1'h0; // @[RA_Mul.scala 417:19:@499.4]
  assign io_matrix_o_1_28 = FA_17_io_cout; // @[RA_Mul.scala 47:10:@498.4]
  assign io_matrix_o_1_29 = 1'h0; // @[RA_Mul.scala 417:19:@504.4]
  assign io_matrix_o_1_30 = 1'h0; // @[RA_Mul.scala 417:19:@514.4]
  assign io_matrix_o_1_31 = FA_18_io_cout; // @[RA_Mul.scala 47:10:@513.4]
  assign io_matrix_o_2_0 = 1'h0; // @[RA_Mul.scala 417:19:@305.4]
  assign io_matrix_o_2_1 = 1'h0; // @[RA_Mul.scala 417:19:@308.4]
  assign io_matrix_o_2_2 = 1'h0; // @[RA_Mul.scala 417:19:@317.4]
  assign io_matrix_o_2_3 = 1'h0; // @[RA_Mul.scala 417:19:@319.4]
  assign io_matrix_o_2_4 = 1'h0; // @[RA_Mul.scala 417:19:@329.4]
  assign io_matrix_o_2_5 = io_matrix_i_1_5; // @[RA_Mul.scala 437:21:@331.4]
  assign io_matrix_o_2_6 = 1'h0; // @[RA_Mul.scala 417:19:@334.4]
  assign io_matrix_o_2_7 = 1'h0; // @[RA_Mul.scala 417:19:@337.4]
  assign io_matrix_o_2_8 = 1'h0; // @[RA_Mul.scala 417:19:@340.4]
  assign io_matrix_o_2_9 = 1'h0; // @[RA_Mul.scala 417:19:@350.4]
  assign io_matrix_o_2_10 = 1'h0; // @[RA_Mul.scala 417:19:@359.4]
  assign io_matrix_o_2_11 = 1'h0; // @[RA_Mul.scala 417:19:@368.4]
  assign io_matrix_o_2_12 = 1'h0; // @[RA_Mul.scala 417:19:@377.4]
  assign io_matrix_o_2_13 = io_matrix_i_3_13; // @[RA_Mul.scala 456:23:@386.4]
  assign io_matrix_o_2_14 = io_matrix_i_3_14; // @[RA_Mul.scala 456:23:@395.4]
  assign io_matrix_o_2_15 = io_matrix_i_3_15; // @[RA_Mul.scala 456:23:@404.4]
  assign io_matrix_o_2_16 = io_matrix_i_3_16; // @[RA_Mul.scala 456:23:@413.4]
  assign io_matrix_o_2_17 = io_matrix_i_3_17; // @[RA_Mul.scala 456:23:@422.4]
  assign io_matrix_o_2_18 = io_matrix_i_3_18; // @[RA_Mul.scala 456:23:@431.4]
  assign io_matrix_o_2_19 = io_matrix_i_3_19; // @[RA_Mul.scala 456:23:@440.4]
  assign io_matrix_o_2_20 = io_matrix_i_3_20; // @[RA_Mul.scala 456:23:@449.4]
  assign io_matrix_o_2_21 = io_matrix_i_3_21; // @[RA_Mul.scala 456:23:@458.4]
  assign io_matrix_o_2_22 = 1'h0; // @[RA_Mul.scala 417:19:@467.4]
  assign io_matrix_o_2_23 = io_matrix_i_3_23; // @[RA_Mul.scala 463:22:@476.4]
  assign io_matrix_o_2_24 = 1'h0; // @[RA_Mul.scala 417:19:@485.4]
  assign io_matrix_o_2_25 = io_matrix_i_1_25; // @[RA_Mul.scala 469:22:@487.4]
  assign io_matrix_o_2_26 = 1'h0; // @[RA_Mul.scala 417:19:@490.4]
  assign io_matrix_o_2_27 = 1'h0; // @[RA_Mul.scala 417:19:@500.4]
  assign io_matrix_o_2_28 = io_matrix_i_1_28; // @[RA_Mul.scala 479:22:@502.4]
  assign io_matrix_o_2_29 = 1'h0; // @[RA_Mul.scala 417:19:@505.4]
  assign io_matrix_o_2_30 = 1'h0; // @[RA_Mul.scala 417:19:@515.4]
  assign io_matrix_o_2_31 = 1'h0; // @[RA_Mul.scala 417:19:@517.4]
  assign HA_io_a = io_matrix_i_0_2; // @[RA_Mul.scala 19:14:@312.4]
  assign HA_io_b = io_matrix_i_1_2; // @[RA_Mul.scala 20:14:@313.4]
  assign FA_io_a = io_matrix_i_0_4; // @[RA_Mul.scala 43:14:@323.4]
  assign FA_io_b = io_matrix_i_1_4; // @[RA_Mul.scala 44:14:@324.4]
  assign FA_io_cin = io_matrix_i_2_4; // @[RA_Mul.scala 45:16:@325.4]
  assign FA_1_io_a = io_matrix_i_0_9; // @[RA_Mul.scala 43:14:@344.4]
  assign FA_1_io_b = io_matrix_i_1_9; // @[RA_Mul.scala 44:14:@345.4]
  assign FA_1_io_cin = io_matrix_i_2_9; // @[RA_Mul.scala 45:16:@346.4]
  assign FA_2_io_a = io_matrix_i_0_10; // @[RA_Mul.scala 43:14:@354.4]
  assign FA_2_io_b = io_matrix_i_1_10; // @[RA_Mul.scala 44:14:@355.4]
  assign FA_2_io_cin = io_matrix_i_2_10; // @[RA_Mul.scala 45:16:@356.4]
  assign FA_3_io_a = io_matrix_i_0_11; // @[RA_Mul.scala 43:14:@363.4]
  assign FA_3_io_b = io_matrix_i_1_11; // @[RA_Mul.scala 44:14:@364.4]
  assign FA_3_io_cin = io_matrix_i_2_11; // @[RA_Mul.scala 45:16:@365.4]
  assign FA_4_io_a = io_matrix_i_0_12; // @[RA_Mul.scala 43:14:@372.4]
  assign FA_4_io_b = io_matrix_i_1_12; // @[RA_Mul.scala 44:14:@373.4]
  assign FA_4_io_cin = io_matrix_i_2_12; // @[RA_Mul.scala 45:16:@374.4]
  assign FA_5_io_a = io_matrix_i_0_13; // @[RA_Mul.scala 43:14:@381.4]
  assign FA_5_io_b = io_matrix_i_1_13; // @[RA_Mul.scala 44:14:@382.4]
  assign FA_5_io_cin = io_matrix_i_2_13; // @[RA_Mul.scala 45:16:@383.4]
  assign FA_6_io_a = io_matrix_i_0_14; // @[RA_Mul.scala 43:14:@390.4]
  assign FA_6_io_b = io_matrix_i_1_14; // @[RA_Mul.scala 44:14:@391.4]
  assign FA_6_io_cin = io_matrix_i_2_14; // @[RA_Mul.scala 45:16:@392.4]
  assign FA_7_io_a = io_matrix_i_0_15; // @[RA_Mul.scala 43:14:@399.4]
  assign FA_7_io_b = io_matrix_i_1_15; // @[RA_Mul.scala 44:14:@400.4]
  assign FA_7_io_cin = io_matrix_i_2_15; // @[RA_Mul.scala 45:16:@401.4]
  assign FA_8_io_a = io_matrix_i_0_16; // @[RA_Mul.scala 43:14:@408.4]
  assign FA_8_io_b = io_matrix_i_1_16; // @[RA_Mul.scala 44:14:@409.4]
  assign FA_8_io_cin = io_matrix_i_2_16; // @[RA_Mul.scala 45:16:@410.4]
  assign FA_9_io_a = io_matrix_i_0_17; // @[RA_Mul.scala 43:14:@417.4]
  assign FA_9_io_b = io_matrix_i_1_17; // @[RA_Mul.scala 44:14:@418.4]
  assign FA_9_io_cin = io_matrix_i_2_17; // @[RA_Mul.scala 45:16:@419.4]
  assign FA_10_io_a = io_matrix_i_0_18; // @[RA_Mul.scala 43:14:@426.4]
  assign FA_10_io_b = io_matrix_i_1_18; // @[RA_Mul.scala 44:14:@427.4]
  assign FA_10_io_cin = io_matrix_i_2_18; // @[RA_Mul.scala 45:16:@428.4]
  assign FA_11_io_a = io_matrix_i_0_19; // @[RA_Mul.scala 43:14:@435.4]
  assign FA_11_io_b = io_matrix_i_1_19; // @[RA_Mul.scala 44:14:@436.4]
  assign FA_11_io_cin = io_matrix_i_2_19; // @[RA_Mul.scala 45:16:@437.4]
  assign FA_12_io_a = io_matrix_i_0_20; // @[RA_Mul.scala 43:14:@444.4]
  assign FA_12_io_b = io_matrix_i_1_20; // @[RA_Mul.scala 44:14:@445.4]
  assign FA_12_io_cin = io_matrix_i_2_20; // @[RA_Mul.scala 45:16:@446.4]
  assign FA_13_io_a = io_matrix_i_0_21; // @[RA_Mul.scala 43:14:@453.4]
  assign FA_13_io_b = io_matrix_i_1_21; // @[RA_Mul.scala 44:14:@454.4]
  assign FA_13_io_cin = io_matrix_i_2_21; // @[RA_Mul.scala 45:16:@455.4]
  assign FA_14_io_a = io_matrix_i_0_22; // @[RA_Mul.scala 43:14:@462.4]
  assign FA_14_io_b = io_matrix_i_1_22; // @[RA_Mul.scala 44:14:@463.4]
  assign FA_14_io_cin = io_matrix_i_2_22; // @[RA_Mul.scala 45:16:@464.4]
  assign FA_15_io_a = io_matrix_i_0_23; // @[RA_Mul.scala 43:14:@471.4]
  assign FA_15_io_b = io_matrix_i_1_23; // @[RA_Mul.scala 44:14:@472.4]
  assign FA_15_io_cin = io_matrix_i_2_23; // @[RA_Mul.scala 45:16:@473.4]
  assign FA_16_io_a = io_matrix_i_0_24; // @[RA_Mul.scala 43:14:@480.4]
  assign FA_16_io_b = io_matrix_i_1_24; // @[RA_Mul.scala 44:14:@481.4]
  assign FA_16_io_cin = io_matrix_i_2_24; // @[RA_Mul.scala 45:16:@482.4]
  assign FA_17_io_a = io_matrix_i_0_27; // @[RA_Mul.scala 43:14:@494.4]
  assign FA_17_io_b = io_matrix_i_1_27; // @[RA_Mul.scala 44:14:@495.4]
  assign FA_17_io_cin = io_matrix_i_2_27; // @[RA_Mul.scala 45:16:@496.4]
  assign FA_18_io_a = io_matrix_i_0_30; // @[RA_Mul.scala 43:14:@509.4]
  assign FA_18_io_b = io_matrix_i_1_30; // @[RA_Mul.scala 44:14:@510.4]
  assign FA_18_io_cin = io_matrix_i_2_30; // @[RA_Mul.scala 45:16:@511.4]
endmodule
