module BoothEncoder_radix4( // @[:@3.2]
  output [2:0]  io_eB_0, // @[:@6.4]
  output [2:0]  io_eB_1, // @[:@6.4]
  output [2:0]  io_eB_2, // @[:@6.4]
  output [2:0]  io_eB_3, // @[:@6.4]
  output [2:0]  io_eB_4, // @[:@6.4]
  output [2:0]  io_eB_5, // @[:@6.4]
  output [2:0]  io_eB_6, // @[:@6.4]
  output [2:0]  io_eB_7, // @[:@6.4]
  input  [15:0] io_B // @[:@6.4]
);
  wire [16:0] B_ext; // @[Cat.scala 30:58:@8.4]
  wire  _T_34; // @[RA_Mul.scala 69:29:@9.4]
  wire  _T_35; // @[RA_Mul.scala 69:50:@10.4]
  wire  _T_36; // @[RA_Mul.scala 69:69:@11.4]
  wire  _T_37; // @[RA_Mul.scala 69:62:@12.4]
  wire  _T_38; // @[RA_Mul.scala 69:43:@13.4]
  wire  _T_39; // @[RA_Mul.scala 69:41:@14.4]
  wire  _T_42; // @[RA_Mul.scala 70:28:@17.4]
  wire  _T_43; // @[RA_Mul.scala 70:25:@18.4]
  wire  _T_45; // @[RA_Mul.scala 70:50:@20.4]
  wire  _T_46; // @[RA_Mul.scala 70:47:@21.4]
  wire  _T_48; // @[RA_Mul.scala 70:70:@23.4]
  wire  _T_50; // @[RA_Mul.scala 70:89:@25.4]
  wire  _T_52; // @[RA_Mul.scala 70:108:@27.4]
  wire  _T_53; // @[RA_Mul.scala 70:66:@28.4]
  wire  _T_56; // @[RA_Mul.scala 71:24:@31.4]
  wire [1:0] _T_57; // @[Cat.scala 30:58:@32.4]
  wire  _T_59; // @[RA_Mul.scala 69:29:@35.4]
  wire  _T_60; // @[RA_Mul.scala 69:50:@36.4]
  wire  _T_62; // @[RA_Mul.scala 69:62:@38.4]
  wire  _T_63; // @[RA_Mul.scala 69:43:@39.4]
  wire  _T_64; // @[RA_Mul.scala 69:41:@40.4]
  wire  _T_67; // @[RA_Mul.scala 70:28:@43.4]
  wire  _T_68; // @[RA_Mul.scala 70:25:@44.4]
  wire  _T_71; // @[RA_Mul.scala 70:47:@47.4]
  wire  _T_73; // @[RA_Mul.scala 70:70:@49.4]
  wire  _T_75; // @[RA_Mul.scala 70:89:@51.4]
  wire  _T_77; // @[RA_Mul.scala 70:108:@53.4]
  wire  _T_78; // @[RA_Mul.scala 70:66:@54.4]
  wire  _T_81; // @[RA_Mul.scala 71:24:@57.4]
  wire [1:0] _T_82; // @[Cat.scala 30:58:@58.4]
  wire  _T_84; // @[RA_Mul.scala 69:29:@61.4]
  wire  _T_85; // @[RA_Mul.scala 69:50:@62.4]
  wire  _T_87; // @[RA_Mul.scala 69:62:@64.4]
  wire  _T_88; // @[RA_Mul.scala 69:43:@65.4]
  wire  _T_89; // @[RA_Mul.scala 69:41:@66.4]
  wire  _T_92; // @[RA_Mul.scala 70:28:@69.4]
  wire  _T_93; // @[RA_Mul.scala 70:25:@70.4]
  wire  _T_96; // @[RA_Mul.scala 70:47:@73.4]
  wire  _T_98; // @[RA_Mul.scala 70:70:@75.4]
  wire  _T_100; // @[RA_Mul.scala 70:89:@77.4]
  wire  _T_102; // @[RA_Mul.scala 70:108:@79.4]
  wire  _T_103; // @[RA_Mul.scala 70:66:@80.4]
  wire  _T_106; // @[RA_Mul.scala 71:24:@83.4]
  wire [1:0] _T_107; // @[Cat.scala 30:58:@84.4]
  wire  _T_109; // @[RA_Mul.scala 69:29:@87.4]
  wire  _T_110; // @[RA_Mul.scala 69:50:@88.4]
  wire  _T_112; // @[RA_Mul.scala 69:62:@90.4]
  wire  _T_113; // @[RA_Mul.scala 69:43:@91.4]
  wire  _T_114; // @[RA_Mul.scala 69:41:@92.4]
  wire  _T_117; // @[RA_Mul.scala 70:28:@95.4]
  wire  _T_118; // @[RA_Mul.scala 70:25:@96.4]
  wire  _T_121; // @[RA_Mul.scala 70:47:@99.4]
  wire  _T_123; // @[RA_Mul.scala 70:70:@101.4]
  wire  _T_125; // @[RA_Mul.scala 70:89:@103.4]
  wire  _T_127; // @[RA_Mul.scala 70:108:@105.4]
  wire  _T_128; // @[RA_Mul.scala 70:66:@106.4]
  wire  _T_131; // @[RA_Mul.scala 71:24:@109.4]
  wire [1:0] _T_132; // @[Cat.scala 30:58:@110.4]
  wire  _T_134; // @[RA_Mul.scala 69:29:@113.4]
  wire  _T_135; // @[RA_Mul.scala 69:50:@114.4]
  wire  _T_137; // @[RA_Mul.scala 69:62:@116.4]
  wire  _T_138; // @[RA_Mul.scala 69:43:@117.4]
  wire  _T_139; // @[RA_Mul.scala 69:41:@118.4]
  wire  _T_142; // @[RA_Mul.scala 70:28:@121.4]
  wire  _T_143; // @[RA_Mul.scala 70:25:@122.4]
  wire  _T_146; // @[RA_Mul.scala 70:47:@125.4]
  wire  _T_148; // @[RA_Mul.scala 70:70:@127.4]
  wire  _T_150; // @[RA_Mul.scala 70:89:@129.4]
  wire  _T_152; // @[RA_Mul.scala 70:108:@131.4]
  wire  _T_153; // @[RA_Mul.scala 70:66:@132.4]
  wire  _T_156; // @[RA_Mul.scala 71:24:@135.4]
  wire [1:0] _T_157; // @[Cat.scala 30:58:@136.4]
  wire  _T_159; // @[RA_Mul.scala 69:29:@139.4]
  wire  _T_160; // @[RA_Mul.scala 69:50:@140.4]
  wire  _T_162; // @[RA_Mul.scala 69:62:@142.4]
  wire  _T_163; // @[RA_Mul.scala 69:43:@143.4]
  wire  _T_164; // @[RA_Mul.scala 69:41:@144.4]
  wire  _T_167; // @[RA_Mul.scala 70:28:@147.4]
  wire  _T_168; // @[RA_Mul.scala 70:25:@148.4]
  wire  _T_171; // @[RA_Mul.scala 70:47:@151.4]
  wire  _T_173; // @[RA_Mul.scala 70:70:@153.4]
  wire  _T_175; // @[RA_Mul.scala 70:89:@155.4]
  wire  _T_177; // @[RA_Mul.scala 70:108:@157.4]
  wire  _T_178; // @[RA_Mul.scala 70:66:@158.4]
  wire  _T_181; // @[RA_Mul.scala 71:24:@161.4]
  wire [1:0] _T_182; // @[Cat.scala 30:58:@162.4]
  wire  _T_184; // @[RA_Mul.scala 69:29:@165.4]
  wire  _T_185; // @[RA_Mul.scala 69:50:@166.4]
  wire  _T_187; // @[RA_Mul.scala 69:62:@168.4]
  wire  _T_188; // @[RA_Mul.scala 69:43:@169.4]
  wire  _T_189; // @[RA_Mul.scala 69:41:@170.4]
  wire  _T_192; // @[RA_Mul.scala 70:28:@173.4]
  wire  _T_193; // @[RA_Mul.scala 70:25:@174.4]
  wire  _T_196; // @[RA_Mul.scala 70:47:@177.4]
  wire  _T_198; // @[RA_Mul.scala 70:70:@179.4]
  wire  _T_200; // @[RA_Mul.scala 70:89:@181.4]
  wire  _T_202; // @[RA_Mul.scala 70:108:@183.4]
  wire  _T_203; // @[RA_Mul.scala 70:66:@184.4]
  wire  _T_206; // @[RA_Mul.scala 71:24:@187.4]
  wire [1:0] _T_207; // @[Cat.scala 30:58:@188.4]
  wire  _T_209; // @[RA_Mul.scala 69:29:@191.4]
  wire  _T_210; // @[RA_Mul.scala 69:50:@192.4]
  wire  _T_212; // @[RA_Mul.scala 69:62:@194.4]
  wire  _T_213; // @[RA_Mul.scala 69:43:@195.4]
  wire  _T_214; // @[RA_Mul.scala 69:41:@196.4]
  wire  _T_217; // @[RA_Mul.scala 70:28:@199.4]
  wire  _T_218; // @[RA_Mul.scala 70:25:@200.4]
  wire  _T_221; // @[RA_Mul.scala 70:47:@203.4]
  wire  _T_223; // @[RA_Mul.scala 70:70:@205.4]
  wire  _T_225; // @[RA_Mul.scala 70:89:@207.4]
  wire  _T_227; // @[RA_Mul.scala 70:108:@209.4]
  wire  _T_228; // @[RA_Mul.scala 70:66:@210.4]
  wire  _T_231; // @[RA_Mul.scala 71:24:@213.4]
  wire [1:0] _T_232; // @[Cat.scala 30:58:@214.4]
  assign B_ext = {io_B,1'h0}; // @[Cat.scala 30:58:@8.4]
  assign _T_34 = B_ext[2]; // @[RA_Mul.scala 69:29:@9.4]
  assign _T_35 = B_ext[1]; // @[RA_Mul.scala 69:50:@10.4]
  assign _T_36 = B_ext[0]; // @[RA_Mul.scala 69:69:@11.4]
  assign _T_37 = _T_35 & _T_36; // @[RA_Mul.scala 69:62:@12.4]
  assign _T_38 = ~ _T_37; // @[RA_Mul.scala 69:43:@13.4]
  assign _T_39 = _T_34 & _T_38; // @[RA_Mul.scala 69:41:@14.4]
  assign _T_42 = ~ _T_35; // @[RA_Mul.scala 70:28:@17.4]
  assign _T_43 = _T_34 & _T_42; // @[RA_Mul.scala 70:25:@18.4]
  assign _T_45 = ~ _T_36; // @[RA_Mul.scala 70:50:@20.4]
  assign _T_46 = _T_43 & _T_45; // @[RA_Mul.scala 70:47:@21.4]
  assign _T_48 = ~ _T_34; // @[RA_Mul.scala 70:70:@23.4]
  assign _T_50 = _T_48 & _T_35; // @[RA_Mul.scala 70:89:@25.4]
  assign _T_52 = _T_50 & _T_36; // @[RA_Mul.scala 70:108:@27.4]
  assign _T_53 = _T_46 | _T_52; // @[RA_Mul.scala 70:66:@28.4]
  assign _T_56 = _T_35 ^ _T_36; // @[RA_Mul.scala 71:24:@31.4]
  assign _T_57 = {_T_39,_T_53}; // @[Cat.scala 30:58:@32.4]
  assign _T_59 = B_ext[4]; // @[RA_Mul.scala 69:29:@35.4]
  assign _T_60 = B_ext[3]; // @[RA_Mul.scala 69:50:@36.4]
  assign _T_62 = _T_60 & _T_34; // @[RA_Mul.scala 69:62:@38.4]
  assign _T_63 = ~ _T_62; // @[RA_Mul.scala 69:43:@39.4]
  assign _T_64 = _T_59 & _T_63; // @[RA_Mul.scala 69:41:@40.4]
  assign _T_67 = ~ _T_60; // @[RA_Mul.scala 70:28:@43.4]
  assign _T_68 = _T_59 & _T_67; // @[RA_Mul.scala 70:25:@44.4]
  assign _T_71 = _T_68 & _T_48; // @[RA_Mul.scala 70:47:@47.4]
  assign _T_73 = ~ _T_59; // @[RA_Mul.scala 70:70:@49.4]
  assign _T_75 = _T_73 & _T_60; // @[RA_Mul.scala 70:89:@51.4]
  assign _T_77 = _T_75 & _T_34; // @[RA_Mul.scala 70:108:@53.4]
  assign _T_78 = _T_71 | _T_77; // @[RA_Mul.scala 70:66:@54.4]
  assign _T_81 = _T_60 ^ _T_34; // @[RA_Mul.scala 71:24:@57.4]
  assign _T_82 = {_T_64,_T_78}; // @[Cat.scala 30:58:@58.4]
  assign _T_84 = B_ext[6]; // @[RA_Mul.scala 69:29:@61.4]
  assign _T_85 = B_ext[5]; // @[RA_Mul.scala 69:50:@62.4]
  assign _T_87 = _T_85 & _T_59; // @[RA_Mul.scala 69:62:@64.4]
  assign _T_88 = ~ _T_87; // @[RA_Mul.scala 69:43:@65.4]
  assign _T_89 = _T_84 & _T_88; // @[RA_Mul.scala 69:41:@66.4]
  assign _T_92 = ~ _T_85; // @[RA_Mul.scala 70:28:@69.4]
  assign _T_93 = _T_84 & _T_92; // @[RA_Mul.scala 70:25:@70.4]
  assign _T_96 = _T_93 & _T_73; // @[RA_Mul.scala 70:47:@73.4]
  assign _T_98 = ~ _T_84; // @[RA_Mul.scala 70:70:@75.4]
  assign _T_100 = _T_98 & _T_85; // @[RA_Mul.scala 70:89:@77.4]
  assign _T_102 = _T_100 & _T_59; // @[RA_Mul.scala 70:108:@79.4]
  assign _T_103 = _T_96 | _T_102; // @[RA_Mul.scala 70:66:@80.4]
  assign _T_106 = _T_85 ^ _T_59; // @[RA_Mul.scala 71:24:@83.4]
  assign _T_107 = {_T_89,_T_103}; // @[Cat.scala 30:58:@84.4]
  assign _T_109 = B_ext[8]; // @[RA_Mul.scala 69:29:@87.4]
  assign _T_110 = B_ext[7]; // @[RA_Mul.scala 69:50:@88.4]
  assign _T_112 = _T_110 & _T_84; // @[RA_Mul.scala 69:62:@90.4]
  assign _T_113 = ~ _T_112; // @[RA_Mul.scala 69:43:@91.4]
  assign _T_114 = _T_109 & _T_113; // @[RA_Mul.scala 69:41:@92.4]
  assign _T_117 = ~ _T_110; // @[RA_Mul.scala 70:28:@95.4]
  assign _T_118 = _T_109 & _T_117; // @[RA_Mul.scala 70:25:@96.4]
  assign _T_121 = _T_118 & _T_98; // @[RA_Mul.scala 70:47:@99.4]
  assign _T_123 = ~ _T_109; // @[RA_Mul.scala 70:70:@101.4]
  assign _T_125 = _T_123 & _T_110; // @[RA_Mul.scala 70:89:@103.4]
  assign _T_127 = _T_125 & _T_84; // @[RA_Mul.scala 70:108:@105.4]
  assign _T_128 = _T_121 | _T_127; // @[RA_Mul.scala 70:66:@106.4]
  assign _T_131 = _T_110 ^ _T_84; // @[RA_Mul.scala 71:24:@109.4]
  assign _T_132 = {_T_114,_T_128}; // @[Cat.scala 30:58:@110.4]
  assign _T_134 = B_ext[10]; // @[RA_Mul.scala 69:29:@113.4]
  assign _T_135 = B_ext[9]; // @[RA_Mul.scala 69:50:@114.4]
  assign _T_137 = _T_135 & _T_109; // @[RA_Mul.scala 69:62:@116.4]
  assign _T_138 = ~ _T_137; // @[RA_Mul.scala 69:43:@117.4]
  assign _T_139 = _T_134 & _T_138; // @[RA_Mul.scala 69:41:@118.4]
  assign _T_142 = ~ _T_135; // @[RA_Mul.scala 70:28:@121.4]
  assign _T_143 = _T_134 & _T_142; // @[RA_Mul.scala 70:25:@122.4]
  assign _T_146 = _T_143 & _T_123; // @[RA_Mul.scala 70:47:@125.4]
  assign _T_148 = ~ _T_134; // @[RA_Mul.scala 70:70:@127.4]
  assign _T_150 = _T_148 & _T_135; // @[RA_Mul.scala 70:89:@129.4]
  assign _T_152 = _T_150 & _T_109; // @[RA_Mul.scala 70:108:@131.4]
  assign _T_153 = _T_146 | _T_152; // @[RA_Mul.scala 70:66:@132.4]
  assign _T_156 = _T_135 ^ _T_109; // @[RA_Mul.scala 71:24:@135.4]
  assign _T_157 = {_T_139,_T_153}; // @[Cat.scala 30:58:@136.4]
  assign _T_159 = B_ext[12]; // @[RA_Mul.scala 69:29:@139.4]
  assign _T_160 = B_ext[11]; // @[RA_Mul.scala 69:50:@140.4]
  assign _T_162 = _T_160 & _T_134; // @[RA_Mul.scala 69:62:@142.4]
  assign _T_163 = ~ _T_162; // @[RA_Mul.scala 69:43:@143.4]
  assign _T_164 = _T_159 & _T_163; // @[RA_Mul.scala 69:41:@144.4]
  assign _T_167 = ~ _T_160; // @[RA_Mul.scala 70:28:@147.4]
  assign _T_168 = _T_159 & _T_167; // @[RA_Mul.scala 70:25:@148.4]
  assign _T_171 = _T_168 & _T_148; // @[RA_Mul.scala 70:47:@151.4]
  assign _T_173 = ~ _T_159; // @[RA_Mul.scala 70:70:@153.4]
  assign _T_175 = _T_173 & _T_160; // @[RA_Mul.scala 70:89:@155.4]
  assign _T_177 = _T_175 & _T_134; // @[RA_Mul.scala 70:108:@157.4]
  assign _T_178 = _T_171 | _T_177; // @[RA_Mul.scala 70:66:@158.4]
  assign _T_181 = _T_160 ^ _T_134; // @[RA_Mul.scala 71:24:@161.4]
  assign _T_182 = {_T_164,_T_178}; // @[Cat.scala 30:58:@162.4]
  assign _T_184 = B_ext[14]; // @[RA_Mul.scala 69:29:@165.4]
  assign _T_185 = B_ext[13]; // @[RA_Mul.scala 69:50:@166.4]
  assign _T_187 = _T_185 & _T_159; // @[RA_Mul.scala 69:62:@168.4]
  assign _T_188 = ~ _T_187; // @[RA_Mul.scala 69:43:@169.4]
  assign _T_189 = _T_184 & _T_188; // @[RA_Mul.scala 69:41:@170.4]
  assign _T_192 = ~ _T_185; // @[RA_Mul.scala 70:28:@173.4]
  assign _T_193 = _T_184 & _T_192; // @[RA_Mul.scala 70:25:@174.4]
  assign _T_196 = _T_193 & _T_173; // @[RA_Mul.scala 70:47:@177.4]
  assign _T_198 = ~ _T_184; // @[RA_Mul.scala 70:70:@179.4]
  assign _T_200 = _T_198 & _T_185; // @[RA_Mul.scala 70:89:@181.4]
  assign _T_202 = _T_200 & _T_159; // @[RA_Mul.scala 70:108:@183.4]
  assign _T_203 = _T_196 | _T_202; // @[RA_Mul.scala 70:66:@184.4]
  assign _T_206 = _T_185 ^ _T_159; // @[RA_Mul.scala 71:24:@187.4]
  assign _T_207 = {_T_189,_T_203}; // @[Cat.scala 30:58:@188.4]
  assign _T_209 = B_ext[16]; // @[RA_Mul.scala 69:29:@191.4]
  assign _T_210 = B_ext[15]; // @[RA_Mul.scala 69:50:@192.4]
  assign _T_212 = _T_210 & _T_184; // @[RA_Mul.scala 69:62:@194.4]
  assign _T_213 = ~ _T_212; // @[RA_Mul.scala 69:43:@195.4]
  assign _T_214 = _T_209 & _T_213; // @[RA_Mul.scala 69:41:@196.4]
  assign _T_217 = ~ _T_210; // @[RA_Mul.scala 70:28:@199.4]
  assign _T_218 = _T_209 & _T_217; // @[RA_Mul.scala 70:25:@200.4]
  assign _T_221 = _T_218 & _T_198; // @[RA_Mul.scala 70:47:@203.4]
  assign _T_223 = ~ _T_209; // @[RA_Mul.scala 70:70:@205.4]
  assign _T_225 = _T_223 & _T_210; // @[RA_Mul.scala 70:89:@207.4]
  assign _T_227 = _T_225 & _T_184; // @[RA_Mul.scala 70:108:@209.4]
  assign _T_228 = _T_221 | _T_227; // @[RA_Mul.scala 70:66:@210.4]
  assign _T_231 = _T_210 ^ _T_184; // @[RA_Mul.scala 71:24:@213.4]
  assign _T_232 = {_T_214,_T_228}; // @[Cat.scala 30:58:@214.4]
  assign io_eB_0 = {_T_57,_T_56}; // @[RA_Mul.scala 69:14:@34.4]
  assign io_eB_1 = {_T_82,_T_81}; // @[RA_Mul.scala 69:14:@60.4]
  assign io_eB_2 = {_T_107,_T_106}; // @[RA_Mul.scala 69:14:@86.4]
  assign io_eB_3 = {_T_132,_T_131}; // @[RA_Mul.scala 69:14:@112.4]
  assign io_eB_4 = {_T_157,_T_156}; // @[RA_Mul.scala 69:14:@138.4]
  assign io_eB_5 = {_T_182,_T_181}; // @[RA_Mul.scala 69:14:@164.4]
  assign io_eB_6 = {_T_207,_T_206}; // @[RA_Mul.scala 69:14:@190.4]
  assign io_eB_7 = {_T_232,_T_231}; // @[RA_Mul.scala 69:14:@216.4]
endmodule
module PPGen( // @[:@218.2]
  output [15:0] io_PP_0, // @[:@221.4]
  output [15:0] io_PP_1, // @[:@221.4]
  output [15:0] io_PP_2, // @[:@221.4]
  output [15:0] io_PP_3, // @[:@221.4]
  output [15:0] io_PP_4, // @[:@221.4]
  output [15:0] io_PP_5, // @[:@221.4]
  output [15:0] io_PP_6, // @[:@221.4]
  output [15:0] io_PP_7, // @[:@221.4]
  output [7:0]  io_SC, // @[:@221.4]
  output [7:0]  io_S, // @[:@221.4]
  input  [2:0]  io_eB_0, // @[:@221.4]
  input  [2:0]  io_eB_1, // @[:@221.4]
  input  [2:0]  io_eB_2, // @[:@221.4]
  input  [2:0]  io_eB_3, // @[:@221.4]
  input  [2:0]  io_eB_4, // @[:@221.4]
  input  [2:0]  io_eB_5, // @[:@221.4]
  input  [2:0]  io_eB_6, // @[:@221.4]
  input  [2:0]  io_eB_7, // @[:@221.4]
  input  [15:0] io_A // @[:@221.4]
);
  wire  _T_93; // @[RA_Mul.scala 125:19:@226.4]
  wire  _T_95; // @[RA_Mul.scala 125:44:@227.4]
  wire  _T_96; // @[RA_Mul.scala 125:32:@228.4]
  wire  _T_99; // @[RA_Mul.scala 127:25:@233.6]
  wire  _T_101; // @[RA_Mul.scala 129:25:@238.8]
  wire [16:0] _GEN_56; // @[RA_Mul.scala 130:25:@240.10]
  wire [16:0] _T_102; // @[RA_Mul.scala 130:25:@240.10]
  wire [15:0] _T_103; // @[RA_Mul.scala 130:30:@241.10]
  wire  _T_105; // @[RA_Mul.scala 131:25:@245.10]
  wire [15:0] _T_106; // @[RA_Mul.scala 132:19:@247.12]
  wire  _T_108; // @[RA_Mul.scala 133:25:@251.12]
  wire [15:0] _T_111; // @[RA_Mul.scala 134:19:@255.14]
  wire [15:0] _GEN_0; // @[RA_Mul.scala 133:38:@252.12]
  wire [15:0] _GEN_1; // @[RA_Mul.scala 131:39:@246.10]
  wire [15:0] _GEN_2; // @[RA_Mul.scala 129:39:@239.8]
  wire [15:0] _GEN_3; // @[RA_Mul.scala 127:39:@234.6]
  wire  S_v_0; // @[RA_Mul.scala 139:23:@261.4]
  wire  _T_118; // @[RA_Mul.scala 142:41:@265.4]
  wire  _T_119; // @[RA_Mul.scala 142:33:@266.4]
  wire  _T_120; // @[RA_Mul.scala 142:57:@267.4]
  wire  _T_122; // @[RA_Mul.scala 142:67:@268.4]
  wire  _T_123; // @[RA_Mul.scala 142:49:@269.4]
  wire  _T_127; // @[RA_Mul.scala 144:28:@275.6]
  wire  _T_128; // @[RA_Mul.scala 144:48:@276.6]
  wire  _T_129; // @[RA_Mul.scala 144:60:@277.6]
  wire  _T_130; // @[RA_Mul.scala 144:51:@278.6]
  wire  _T_133; // @[RA_Mul.scala 144:36:@280.6]
  wire  _T_137; // @[RA_Mul.scala 144:73:@283.6]
  wire  _GEN_5; // @[RA_Mul.scala 144:98:@284.6]
  wire  SC_v_0; // @[RA_Mul.scala 142:75:@270.4]
  wire  _T_141; // @[RA_Mul.scala 125:19:@290.4]
  wire  _T_143; // @[RA_Mul.scala 125:44:@291.4]
  wire  _T_144; // @[RA_Mul.scala 125:32:@292.4]
  wire  _T_147; // @[RA_Mul.scala 127:25:@297.6]
  wire  _T_149; // @[RA_Mul.scala 129:25:@302.8]
  wire  _T_153; // @[RA_Mul.scala 131:25:@309.10]
  wire  _T_156; // @[RA_Mul.scala 133:25:@315.12]
  wire [15:0] _GEN_7; // @[RA_Mul.scala 133:38:@316.12]
  wire [15:0] _GEN_8; // @[RA_Mul.scala 131:39:@310.10]
  wire [15:0] _GEN_9; // @[RA_Mul.scala 129:39:@303.8]
  wire [15:0] _GEN_10; // @[RA_Mul.scala 127:39:@298.6]
  wire  S_v_1; // @[RA_Mul.scala 139:23:@325.4]
  wire  _T_167; // @[RA_Mul.scala 142:33:@330.4]
  wire  _T_171; // @[RA_Mul.scala 142:49:@333.4]
  wire  _T_175; // @[RA_Mul.scala 144:28:@339.6]
  wire  _T_176; // @[RA_Mul.scala 144:48:@340.6]
  wire  _T_177; // @[RA_Mul.scala 144:60:@341.6]
  wire  _T_178; // @[RA_Mul.scala 144:51:@342.6]
  wire  _T_181; // @[RA_Mul.scala 144:36:@344.6]
  wire  _T_185; // @[RA_Mul.scala 144:73:@347.6]
  wire  _GEN_12; // @[RA_Mul.scala 144:98:@348.6]
  wire  SC_v_1; // @[RA_Mul.scala 142:75:@334.4]
  wire  _T_189; // @[RA_Mul.scala 125:19:@354.4]
  wire  _T_191; // @[RA_Mul.scala 125:44:@355.4]
  wire  _T_192; // @[RA_Mul.scala 125:32:@356.4]
  wire  _T_195; // @[RA_Mul.scala 127:25:@361.6]
  wire  _T_197; // @[RA_Mul.scala 129:25:@366.8]
  wire  _T_201; // @[RA_Mul.scala 131:25:@373.10]
  wire  _T_204; // @[RA_Mul.scala 133:25:@379.12]
  wire [15:0] _GEN_14; // @[RA_Mul.scala 133:38:@380.12]
  wire [15:0] _GEN_15; // @[RA_Mul.scala 131:39:@374.10]
  wire [15:0] _GEN_16; // @[RA_Mul.scala 129:39:@367.8]
  wire [15:0] _GEN_17; // @[RA_Mul.scala 127:39:@362.6]
  wire  S_v_2; // @[RA_Mul.scala 139:23:@389.4]
  wire  _T_215; // @[RA_Mul.scala 142:33:@394.4]
  wire  _T_219; // @[RA_Mul.scala 142:49:@397.4]
  wire  _T_223; // @[RA_Mul.scala 144:28:@403.6]
  wire  _T_224; // @[RA_Mul.scala 144:48:@404.6]
  wire  _T_225; // @[RA_Mul.scala 144:60:@405.6]
  wire  _T_226; // @[RA_Mul.scala 144:51:@406.6]
  wire  _T_229; // @[RA_Mul.scala 144:36:@408.6]
  wire  _T_233; // @[RA_Mul.scala 144:73:@411.6]
  wire  _GEN_19; // @[RA_Mul.scala 144:98:@412.6]
  wire  SC_v_2; // @[RA_Mul.scala 142:75:@398.4]
  wire  _T_237; // @[RA_Mul.scala 125:19:@418.4]
  wire  _T_239; // @[RA_Mul.scala 125:44:@419.4]
  wire  _T_240; // @[RA_Mul.scala 125:32:@420.4]
  wire  _T_243; // @[RA_Mul.scala 127:25:@425.6]
  wire  _T_245; // @[RA_Mul.scala 129:25:@430.8]
  wire  _T_249; // @[RA_Mul.scala 131:25:@437.10]
  wire  _T_252; // @[RA_Mul.scala 133:25:@443.12]
  wire [15:0] _GEN_21; // @[RA_Mul.scala 133:38:@444.12]
  wire [15:0] _GEN_22; // @[RA_Mul.scala 131:39:@438.10]
  wire [15:0] _GEN_23; // @[RA_Mul.scala 129:39:@431.8]
  wire [15:0] _GEN_24; // @[RA_Mul.scala 127:39:@426.6]
  wire  S_v_3; // @[RA_Mul.scala 139:23:@453.4]
  wire  _T_263; // @[RA_Mul.scala 142:33:@458.4]
  wire  _T_267; // @[RA_Mul.scala 142:49:@461.4]
  wire  _T_271; // @[RA_Mul.scala 144:28:@467.6]
  wire  _T_272; // @[RA_Mul.scala 144:48:@468.6]
  wire  _T_273; // @[RA_Mul.scala 144:60:@469.6]
  wire  _T_274; // @[RA_Mul.scala 144:51:@470.6]
  wire  _T_277; // @[RA_Mul.scala 144:36:@472.6]
  wire  _T_281; // @[RA_Mul.scala 144:73:@475.6]
  wire  _GEN_26; // @[RA_Mul.scala 144:98:@476.6]
  wire  SC_v_3; // @[RA_Mul.scala 142:75:@462.4]
  wire  _T_285; // @[RA_Mul.scala 125:19:@482.4]
  wire  _T_287; // @[RA_Mul.scala 125:44:@483.4]
  wire  _T_288; // @[RA_Mul.scala 125:32:@484.4]
  wire  _T_291; // @[RA_Mul.scala 127:25:@489.6]
  wire  _T_293; // @[RA_Mul.scala 129:25:@494.8]
  wire  _T_297; // @[RA_Mul.scala 131:25:@501.10]
  wire  _T_300; // @[RA_Mul.scala 133:25:@507.12]
  wire [15:0] _GEN_28; // @[RA_Mul.scala 133:38:@508.12]
  wire [15:0] _GEN_29; // @[RA_Mul.scala 131:39:@502.10]
  wire [15:0] _GEN_30; // @[RA_Mul.scala 129:39:@495.8]
  wire [15:0] _GEN_31; // @[RA_Mul.scala 127:39:@490.6]
  wire  S_v_4; // @[RA_Mul.scala 139:23:@517.4]
  wire  _T_311; // @[RA_Mul.scala 142:33:@522.4]
  wire  _T_315; // @[RA_Mul.scala 142:49:@525.4]
  wire  _T_319; // @[RA_Mul.scala 144:28:@531.6]
  wire  _T_320; // @[RA_Mul.scala 144:48:@532.6]
  wire  _T_321; // @[RA_Mul.scala 144:60:@533.6]
  wire  _T_322; // @[RA_Mul.scala 144:51:@534.6]
  wire  _T_325; // @[RA_Mul.scala 144:36:@536.6]
  wire  _T_329; // @[RA_Mul.scala 144:73:@539.6]
  wire  _GEN_33; // @[RA_Mul.scala 144:98:@540.6]
  wire  SC_v_4; // @[RA_Mul.scala 142:75:@526.4]
  wire  _T_333; // @[RA_Mul.scala 125:19:@546.4]
  wire  _T_335; // @[RA_Mul.scala 125:44:@547.4]
  wire  _T_336; // @[RA_Mul.scala 125:32:@548.4]
  wire  _T_339; // @[RA_Mul.scala 127:25:@553.6]
  wire  _T_341; // @[RA_Mul.scala 129:25:@558.8]
  wire  _T_345; // @[RA_Mul.scala 131:25:@565.10]
  wire  _T_348; // @[RA_Mul.scala 133:25:@571.12]
  wire [15:0] _GEN_35; // @[RA_Mul.scala 133:38:@572.12]
  wire [15:0] _GEN_36; // @[RA_Mul.scala 131:39:@566.10]
  wire [15:0] _GEN_37; // @[RA_Mul.scala 129:39:@559.8]
  wire [15:0] _GEN_38; // @[RA_Mul.scala 127:39:@554.6]
  wire  S_v_5; // @[RA_Mul.scala 139:23:@581.4]
  wire  _T_359; // @[RA_Mul.scala 142:33:@586.4]
  wire  _T_363; // @[RA_Mul.scala 142:49:@589.4]
  wire  _T_367; // @[RA_Mul.scala 144:28:@595.6]
  wire  _T_368; // @[RA_Mul.scala 144:48:@596.6]
  wire  _T_369; // @[RA_Mul.scala 144:60:@597.6]
  wire  _T_370; // @[RA_Mul.scala 144:51:@598.6]
  wire  _T_373; // @[RA_Mul.scala 144:36:@600.6]
  wire  _T_377; // @[RA_Mul.scala 144:73:@603.6]
  wire  _GEN_40; // @[RA_Mul.scala 144:98:@604.6]
  wire  SC_v_5; // @[RA_Mul.scala 142:75:@590.4]
  wire  _T_381; // @[RA_Mul.scala 125:19:@610.4]
  wire  _T_383; // @[RA_Mul.scala 125:44:@611.4]
  wire  _T_384; // @[RA_Mul.scala 125:32:@612.4]
  wire  _T_387; // @[RA_Mul.scala 127:25:@617.6]
  wire  _T_389; // @[RA_Mul.scala 129:25:@622.8]
  wire  _T_393; // @[RA_Mul.scala 131:25:@629.10]
  wire  _T_396; // @[RA_Mul.scala 133:25:@635.12]
  wire [15:0] _GEN_42; // @[RA_Mul.scala 133:38:@636.12]
  wire [15:0] _GEN_43; // @[RA_Mul.scala 131:39:@630.10]
  wire [15:0] _GEN_44; // @[RA_Mul.scala 129:39:@623.8]
  wire [15:0] _GEN_45; // @[RA_Mul.scala 127:39:@618.6]
  wire  S_v_6; // @[RA_Mul.scala 139:23:@645.4]
  wire  _T_407; // @[RA_Mul.scala 142:33:@650.4]
  wire  _T_411; // @[RA_Mul.scala 142:49:@653.4]
  wire  _T_415; // @[RA_Mul.scala 144:28:@659.6]
  wire  _T_416; // @[RA_Mul.scala 144:48:@660.6]
  wire  _T_417; // @[RA_Mul.scala 144:60:@661.6]
  wire  _T_418; // @[RA_Mul.scala 144:51:@662.6]
  wire  _T_421; // @[RA_Mul.scala 144:36:@664.6]
  wire  _T_425; // @[RA_Mul.scala 144:73:@667.6]
  wire  _GEN_47; // @[RA_Mul.scala 144:98:@668.6]
  wire  SC_v_6; // @[RA_Mul.scala 142:75:@654.4]
  wire  _T_429; // @[RA_Mul.scala 125:19:@674.4]
  wire  _T_431; // @[RA_Mul.scala 125:44:@675.4]
  wire  _T_432; // @[RA_Mul.scala 125:32:@676.4]
  wire  _T_435; // @[RA_Mul.scala 127:25:@681.6]
  wire  _T_437; // @[RA_Mul.scala 129:25:@686.8]
  wire  _T_441; // @[RA_Mul.scala 131:25:@693.10]
  wire  _T_444; // @[RA_Mul.scala 133:25:@699.12]
  wire [15:0] _GEN_49; // @[RA_Mul.scala 133:38:@700.12]
  wire [15:0] _GEN_50; // @[RA_Mul.scala 131:39:@694.10]
  wire [15:0] _GEN_51; // @[RA_Mul.scala 129:39:@687.8]
  wire [15:0] _GEN_52; // @[RA_Mul.scala 127:39:@682.6]
  wire  S_v_7; // @[RA_Mul.scala 139:23:@709.4]
  wire  _T_455; // @[RA_Mul.scala 142:33:@714.4]
  wire  _T_459; // @[RA_Mul.scala 142:49:@717.4]
  wire  _T_463; // @[RA_Mul.scala 144:28:@723.6]
  wire  _T_464; // @[RA_Mul.scala 144:48:@724.6]
  wire  _T_465; // @[RA_Mul.scala 144:60:@725.6]
  wire  _T_466; // @[RA_Mul.scala 144:51:@726.6]
  wire  _T_469; // @[RA_Mul.scala 144:36:@728.6]
  wire  _T_473; // @[RA_Mul.scala 144:73:@731.6]
  wire  _GEN_54; // @[RA_Mul.scala 144:98:@732.6]
  wire  SC_v_7; // @[RA_Mul.scala 142:75:@718.4]
  wire [1:0] _T_476; // @[RA_Mul.scala 150:21:@738.4]
  wire [1:0] _T_477; // @[RA_Mul.scala 150:21:@739.4]
  wire [3:0] _T_478; // @[RA_Mul.scala 150:21:@740.4]
  wire [1:0] _T_479; // @[RA_Mul.scala 150:21:@741.4]
  wire [1:0] _T_480; // @[RA_Mul.scala 150:21:@742.4]
  wire [3:0] _T_481; // @[RA_Mul.scala 150:21:@743.4]
  wire [1:0] _T_483; // @[RA_Mul.scala 151:23:@746.4]
  wire [1:0] _T_484; // @[RA_Mul.scala 151:23:@747.4]
  wire [3:0] _T_485; // @[RA_Mul.scala 151:23:@748.4]
  wire [1:0] _T_486; // @[RA_Mul.scala 151:23:@749.4]
  wire [1:0] _T_487; // @[RA_Mul.scala 151:23:@750.4]
  wire [3:0] _T_488; // @[RA_Mul.scala 151:23:@751.4]
  assign _T_93 = io_eB_0 == 3'h0; // @[RA_Mul.scala 125:19:@226.4]
  assign _T_95 = io_eB_0 == 3'h4; // @[RA_Mul.scala 125:44:@227.4]
  assign _T_96 = _T_93 | _T_95; // @[RA_Mul.scala 125:32:@228.4]
  assign _T_99 = io_eB_0 == 3'h1; // @[RA_Mul.scala 127:25:@233.6]
  assign _T_101 = io_eB_0 == 3'h2; // @[RA_Mul.scala 129:25:@238.8]
  assign _GEN_56 = {{1'd0}, io_A}; // @[RA_Mul.scala 130:25:@240.10]
  assign _T_102 = _GEN_56 << 1; // @[RA_Mul.scala 130:25:@240.10]
  assign _T_103 = _T_102[15:0]; // @[RA_Mul.scala 130:30:@241.10]
  assign _T_105 = io_eB_0 == 3'h5; // @[RA_Mul.scala 131:25:@245.10]
  assign _T_106 = ~ io_A; // @[RA_Mul.scala 132:19:@247.12]
  assign _T_108 = io_eB_0 == 3'h6; // @[RA_Mul.scala 133:25:@251.12]
  assign _T_111 = ~ _T_103; // @[RA_Mul.scala 134:19:@255.14]
  assign _GEN_0 = _T_108 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@252.12]
  assign _GEN_1 = _T_105 ? _T_106 : _GEN_0; // @[RA_Mul.scala 131:39:@246.10]
  assign _GEN_2 = _T_101 ? _T_103 : _GEN_1; // @[RA_Mul.scala 129:39:@239.8]
  assign _GEN_3 = _T_99 ? io_A : _GEN_2; // @[RA_Mul.scala 127:39:@234.6]
  assign S_v_0 = io_eB_0[2]; // @[RA_Mul.scala 139:23:@261.4]
  assign _T_118 = io_A != 16'h0; // @[RA_Mul.scala 142:41:@265.4]
  assign _T_119 = S_v_0 & _T_118; // @[RA_Mul.scala 142:33:@266.4]
  assign _T_120 = io_A[15]; // @[RA_Mul.scala 142:57:@267.4]
  assign _T_122 = _T_120 == 1'h0; // @[RA_Mul.scala 142:67:@268.4]
  assign _T_123 = _T_119 & _T_122; // @[RA_Mul.scala 142:49:@269.4]
  assign _T_127 = S_v_0 == 1'h0; // @[RA_Mul.scala 144:28:@275.6]
  assign _T_128 = io_eB_0[1]; // @[RA_Mul.scala 144:48:@276.6]
  assign _T_129 = io_eB_0[0]; // @[RA_Mul.scala 144:60:@277.6]
  assign _T_130 = _T_128 | _T_129; // @[RA_Mul.scala 144:51:@278.6]
  assign _T_133 = _T_127 & _T_130; // @[RA_Mul.scala 144:36:@280.6]
  assign _T_137 = _T_133 & _T_120; // @[RA_Mul.scala 144:73:@283.6]
  assign _GEN_5 = _T_137 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@284.6]
  assign SC_v_0 = _T_123 ? 1'h0 : _GEN_5; // @[RA_Mul.scala 142:75:@270.4]
  assign _T_141 = io_eB_1 == 3'h0; // @[RA_Mul.scala 125:19:@290.4]
  assign _T_143 = io_eB_1 == 3'h4; // @[RA_Mul.scala 125:44:@291.4]
  assign _T_144 = _T_141 | _T_143; // @[RA_Mul.scala 125:32:@292.4]
  assign _T_147 = io_eB_1 == 3'h1; // @[RA_Mul.scala 127:25:@297.6]
  assign _T_149 = io_eB_1 == 3'h2; // @[RA_Mul.scala 129:25:@302.8]
  assign _T_153 = io_eB_1 == 3'h5; // @[RA_Mul.scala 131:25:@309.10]
  assign _T_156 = io_eB_1 == 3'h6; // @[RA_Mul.scala 133:25:@315.12]
  assign _GEN_7 = _T_156 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@316.12]
  assign _GEN_8 = _T_153 ? _T_106 : _GEN_7; // @[RA_Mul.scala 131:39:@310.10]
  assign _GEN_9 = _T_149 ? _T_103 : _GEN_8; // @[RA_Mul.scala 129:39:@303.8]
  assign _GEN_10 = _T_147 ? io_A : _GEN_9; // @[RA_Mul.scala 127:39:@298.6]
  assign S_v_1 = io_eB_1[2]; // @[RA_Mul.scala 139:23:@325.4]
  assign _T_167 = S_v_1 & _T_118; // @[RA_Mul.scala 142:33:@330.4]
  assign _T_171 = _T_167 & _T_122; // @[RA_Mul.scala 142:49:@333.4]
  assign _T_175 = S_v_1 == 1'h0; // @[RA_Mul.scala 144:28:@339.6]
  assign _T_176 = io_eB_1[1]; // @[RA_Mul.scala 144:48:@340.6]
  assign _T_177 = io_eB_1[0]; // @[RA_Mul.scala 144:60:@341.6]
  assign _T_178 = _T_176 | _T_177; // @[RA_Mul.scala 144:51:@342.6]
  assign _T_181 = _T_175 & _T_178; // @[RA_Mul.scala 144:36:@344.6]
  assign _T_185 = _T_181 & _T_120; // @[RA_Mul.scala 144:73:@347.6]
  assign _GEN_12 = _T_185 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@348.6]
  assign SC_v_1 = _T_171 ? 1'h0 : _GEN_12; // @[RA_Mul.scala 142:75:@334.4]
  assign _T_189 = io_eB_2 == 3'h0; // @[RA_Mul.scala 125:19:@354.4]
  assign _T_191 = io_eB_2 == 3'h4; // @[RA_Mul.scala 125:44:@355.4]
  assign _T_192 = _T_189 | _T_191; // @[RA_Mul.scala 125:32:@356.4]
  assign _T_195 = io_eB_2 == 3'h1; // @[RA_Mul.scala 127:25:@361.6]
  assign _T_197 = io_eB_2 == 3'h2; // @[RA_Mul.scala 129:25:@366.8]
  assign _T_201 = io_eB_2 == 3'h5; // @[RA_Mul.scala 131:25:@373.10]
  assign _T_204 = io_eB_2 == 3'h6; // @[RA_Mul.scala 133:25:@379.12]
  assign _GEN_14 = _T_204 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@380.12]
  assign _GEN_15 = _T_201 ? _T_106 : _GEN_14; // @[RA_Mul.scala 131:39:@374.10]
  assign _GEN_16 = _T_197 ? _T_103 : _GEN_15; // @[RA_Mul.scala 129:39:@367.8]
  assign _GEN_17 = _T_195 ? io_A : _GEN_16; // @[RA_Mul.scala 127:39:@362.6]
  assign S_v_2 = io_eB_2[2]; // @[RA_Mul.scala 139:23:@389.4]
  assign _T_215 = S_v_2 & _T_118; // @[RA_Mul.scala 142:33:@394.4]
  assign _T_219 = _T_215 & _T_122; // @[RA_Mul.scala 142:49:@397.4]
  assign _T_223 = S_v_2 == 1'h0; // @[RA_Mul.scala 144:28:@403.6]
  assign _T_224 = io_eB_2[1]; // @[RA_Mul.scala 144:48:@404.6]
  assign _T_225 = io_eB_2[0]; // @[RA_Mul.scala 144:60:@405.6]
  assign _T_226 = _T_224 | _T_225; // @[RA_Mul.scala 144:51:@406.6]
  assign _T_229 = _T_223 & _T_226; // @[RA_Mul.scala 144:36:@408.6]
  assign _T_233 = _T_229 & _T_120; // @[RA_Mul.scala 144:73:@411.6]
  assign _GEN_19 = _T_233 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@412.6]
  assign SC_v_2 = _T_219 ? 1'h0 : _GEN_19; // @[RA_Mul.scala 142:75:@398.4]
  assign _T_237 = io_eB_3 == 3'h0; // @[RA_Mul.scala 125:19:@418.4]
  assign _T_239 = io_eB_3 == 3'h4; // @[RA_Mul.scala 125:44:@419.4]
  assign _T_240 = _T_237 | _T_239; // @[RA_Mul.scala 125:32:@420.4]
  assign _T_243 = io_eB_3 == 3'h1; // @[RA_Mul.scala 127:25:@425.6]
  assign _T_245 = io_eB_3 == 3'h2; // @[RA_Mul.scala 129:25:@430.8]
  assign _T_249 = io_eB_3 == 3'h5; // @[RA_Mul.scala 131:25:@437.10]
  assign _T_252 = io_eB_3 == 3'h6; // @[RA_Mul.scala 133:25:@443.12]
  assign _GEN_21 = _T_252 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@444.12]
  assign _GEN_22 = _T_249 ? _T_106 : _GEN_21; // @[RA_Mul.scala 131:39:@438.10]
  assign _GEN_23 = _T_245 ? _T_103 : _GEN_22; // @[RA_Mul.scala 129:39:@431.8]
  assign _GEN_24 = _T_243 ? io_A : _GEN_23; // @[RA_Mul.scala 127:39:@426.6]
  assign S_v_3 = io_eB_3[2]; // @[RA_Mul.scala 139:23:@453.4]
  assign _T_263 = S_v_3 & _T_118; // @[RA_Mul.scala 142:33:@458.4]
  assign _T_267 = _T_263 & _T_122; // @[RA_Mul.scala 142:49:@461.4]
  assign _T_271 = S_v_3 == 1'h0; // @[RA_Mul.scala 144:28:@467.6]
  assign _T_272 = io_eB_3[1]; // @[RA_Mul.scala 144:48:@468.6]
  assign _T_273 = io_eB_3[0]; // @[RA_Mul.scala 144:60:@469.6]
  assign _T_274 = _T_272 | _T_273; // @[RA_Mul.scala 144:51:@470.6]
  assign _T_277 = _T_271 & _T_274; // @[RA_Mul.scala 144:36:@472.6]
  assign _T_281 = _T_277 & _T_120; // @[RA_Mul.scala 144:73:@475.6]
  assign _GEN_26 = _T_281 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@476.6]
  assign SC_v_3 = _T_267 ? 1'h0 : _GEN_26; // @[RA_Mul.scala 142:75:@462.4]
  assign _T_285 = io_eB_4 == 3'h0; // @[RA_Mul.scala 125:19:@482.4]
  assign _T_287 = io_eB_4 == 3'h4; // @[RA_Mul.scala 125:44:@483.4]
  assign _T_288 = _T_285 | _T_287; // @[RA_Mul.scala 125:32:@484.4]
  assign _T_291 = io_eB_4 == 3'h1; // @[RA_Mul.scala 127:25:@489.6]
  assign _T_293 = io_eB_4 == 3'h2; // @[RA_Mul.scala 129:25:@494.8]
  assign _T_297 = io_eB_4 == 3'h5; // @[RA_Mul.scala 131:25:@501.10]
  assign _T_300 = io_eB_4 == 3'h6; // @[RA_Mul.scala 133:25:@507.12]
  assign _GEN_28 = _T_300 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@508.12]
  assign _GEN_29 = _T_297 ? _T_106 : _GEN_28; // @[RA_Mul.scala 131:39:@502.10]
  assign _GEN_30 = _T_293 ? _T_103 : _GEN_29; // @[RA_Mul.scala 129:39:@495.8]
  assign _GEN_31 = _T_291 ? io_A : _GEN_30; // @[RA_Mul.scala 127:39:@490.6]
  assign S_v_4 = io_eB_4[2]; // @[RA_Mul.scala 139:23:@517.4]
  assign _T_311 = S_v_4 & _T_118; // @[RA_Mul.scala 142:33:@522.4]
  assign _T_315 = _T_311 & _T_122; // @[RA_Mul.scala 142:49:@525.4]
  assign _T_319 = S_v_4 == 1'h0; // @[RA_Mul.scala 144:28:@531.6]
  assign _T_320 = io_eB_4[1]; // @[RA_Mul.scala 144:48:@532.6]
  assign _T_321 = io_eB_4[0]; // @[RA_Mul.scala 144:60:@533.6]
  assign _T_322 = _T_320 | _T_321; // @[RA_Mul.scala 144:51:@534.6]
  assign _T_325 = _T_319 & _T_322; // @[RA_Mul.scala 144:36:@536.6]
  assign _T_329 = _T_325 & _T_120; // @[RA_Mul.scala 144:73:@539.6]
  assign _GEN_33 = _T_329 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@540.6]
  assign SC_v_4 = _T_315 ? 1'h0 : _GEN_33; // @[RA_Mul.scala 142:75:@526.4]
  assign _T_333 = io_eB_5 == 3'h0; // @[RA_Mul.scala 125:19:@546.4]
  assign _T_335 = io_eB_5 == 3'h4; // @[RA_Mul.scala 125:44:@547.4]
  assign _T_336 = _T_333 | _T_335; // @[RA_Mul.scala 125:32:@548.4]
  assign _T_339 = io_eB_5 == 3'h1; // @[RA_Mul.scala 127:25:@553.6]
  assign _T_341 = io_eB_5 == 3'h2; // @[RA_Mul.scala 129:25:@558.8]
  assign _T_345 = io_eB_5 == 3'h5; // @[RA_Mul.scala 131:25:@565.10]
  assign _T_348 = io_eB_5 == 3'h6; // @[RA_Mul.scala 133:25:@571.12]
  assign _GEN_35 = _T_348 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@572.12]
  assign _GEN_36 = _T_345 ? _T_106 : _GEN_35; // @[RA_Mul.scala 131:39:@566.10]
  assign _GEN_37 = _T_341 ? _T_103 : _GEN_36; // @[RA_Mul.scala 129:39:@559.8]
  assign _GEN_38 = _T_339 ? io_A : _GEN_37; // @[RA_Mul.scala 127:39:@554.6]
  assign S_v_5 = io_eB_5[2]; // @[RA_Mul.scala 139:23:@581.4]
  assign _T_359 = S_v_5 & _T_118; // @[RA_Mul.scala 142:33:@586.4]
  assign _T_363 = _T_359 & _T_122; // @[RA_Mul.scala 142:49:@589.4]
  assign _T_367 = S_v_5 == 1'h0; // @[RA_Mul.scala 144:28:@595.6]
  assign _T_368 = io_eB_5[1]; // @[RA_Mul.scala 144:48:@596.6]
  assign _T_369 = io_eB_5[0]; // @[RA_Mul.scala 144:60:@597.6]
  assign _T_370 = _T_368 | _T_369; // @[RA_Mul.scala 144:51:@598.6]
  assign _T_373 = _T_367 & _T_370; // @[RA_Mul.scala 144:36:@600.6]
  assign _T_377 = _T_373 & _T_120; // @[RA_Mul.scala 144:73:@603.6]
  assign _GEN_40 = _T_377 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@604.6]
  assign SC_v_5 = _T_363 ? 1'h0 : _GEN_40; // @[RA_Mul.scala 142:75:@590.4]
  assign _T_381 = io_eB_6 == 3'h0; // @[RA_Mul.scala 125:19:@610.4]
  assign _T_383 = io_eB_6 == 3'h4; // @[RA_Mul.scala 125:44:@611.4]
  assign _T_384 = _T_381 | _T_383; // @[RA_Mul.scala 125:32:@612.4]
  assign _T_387 = io_eB_6 == 3'h1; // @[RA_Mul.scala 127:25:@617.6]
  assign _T_389 = io_eB_6 == 3'h2; // @[RA_Mul.scala 129:25:@622.8]
  assign _T_393 = io_eB_6 == 3'h5; // @[RA_Mul.scala 131:25:@629.10]
  assign _T_396 = io_eB_6 == 3'h6; // @[RA_Mul.scala 133:25:@635.12]
  assign _GEN_42 = _T_396 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@636.12]
  assign _GEN_43 = _T_393 ? _T_106 : _GEN_42; // @[RA_Mul.scala 131:39:@630.10]
  assign _GEN_44 = _T_389 ? _T_103 : _GEN_43; // @[RA_Mul.scala 129:39:@623.8]
  assign _GEN_45 = _T_387 ? io_A : _GEN_44; // @[RA_Mul.scala 127:39:@618.6]
  assign S_v_6 = io_eB_6[2]; // @[RA_Mul.scala 139:23:@645.4]
  assign _T_407 = S_v_6 & _T_118; // @[RA_Mul.scala 142:33:@650.4]
  assign _T_411 = _T_407 & _T_122; // @[RA_Mul.scala 142:49:@653.4]
  assign _T_415 = S_v_6 == 1'h0; // @[RA_Mul.scala 144:28:@659.6]
  assign _T_416 = io_eB_6[1]; // @[RA_Mul.scala 144:48:@660.6]
  assign _T_417 = io_eB_6[0]; // @[RA_Mul.scala 144:60:@661.6]
  assign _T_418 = _T_416 | _T_417; // @[RA_Mul.scala 144:51:@662.6]
  assign _T_421 = _T_415 & _T_418; // @[RA_Mul.scala 144:36:@664.6]
  assign _T_425 = _T_421 & _T_120; // @[RA_Mul.scala 144:73:@667.6]
  assign _GEN_47 = _T_425 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@668.6]
  assign SC_v_6 = _T_411 ? 1'h0 : _GEN_47; // @[RA_Mul.scala 142:75:@654.4]
  assign _T_429 = io_eB_7 == 3'h0; // @[RA_Mul.scala 125:19:@674.4]
  assign _T_431 = io_eB_7 == 3'h4; // @[RA_Mul.scala 125:44:@675.4]
  assign _T_432 = _T_429 | _T_431; // @[RA_Mul.scala 125:32:@676.4]
  assign _T_435 = io_eB_7 == 3'h1; // @[RA_Mul.scala 127:25:@681.6]
  assign _T_437 = io_eB_7 == 3'h2; // @[RA_Mul.scala 129:25:@686.8]
  assign _T_441 = io_eB_7 == 3'h5; // @[RA_Mul.scala 131:25:@693.10]
  assign _T_444 = io_eB_7 == 3'h6; // @[RA_Mul.scala 133:25:@699.12]
  assign _GEN_49 = _T_444 ? _T_111 : 16'h0; // @[RA_Mul.scala 133:38:@700.12]
  assign _GEN_50 = _T_441 ? _T_106 : _GEN_49; // @[RA_Mul.scala 131:39:@694.10]
  assign _GEN_51 = _T_437 ? _T_103 : _GEN_50; // @[RA_Mul.scala 129:39:@687.8]
  assign _GEN_52 = _T_435 ? io_A : _GEN_51; // @[RA_Mul.scala 127:39:@682.6]
  assign S_v_7 = io_eB_7[2]; // @[RA_Mul.scala 139:23:@709.4]
  assign _T_455 = S_v_7 & _T_118; // @[RA_Mul.scala 142:33:@714.4]
  assign _T_459 = _T_455 & _T_122; // @[RA_Mul.scala 142:49:@717.4]
  assign _T_463 = S_v_7 == 1'h0; // @[RA_Mul.scala 144:28:@723.6]
  assign _T_464 = io_eB_7[1]; // @[RA_Mul.scala 144:48:@724.6]
  assign _T_465 = io_eB_7[0]; // @[RA_Mul.scala 144:60:@725.6]
  assign _T_466 = _T_464 | _T_465; // @[RA_Mul.scala 144:51:@726.6]
  assign _T_469 = _T_463 & _T_466; // @[RA_Mul.scala 144:36:@728.6]
  assign _T_473 = _T_469 & _T_120; // @[RA_Mul.scala 144:73:@731.6]
  assign _GEN_54 = _T_473 ? 1'h0 : 1'h1; // @[RA_Mul.scala 144:98:@732.6]
  assign SC_v_7 = _T_459 ? 1'h0 : _GEN_54; // @[RA_Mul.scala 142:75:@718.4]
  assign _T_476 = {S_v_1,S_v_0}; // @[RA_Mul.scala 150:21:@738.4]
  assign _T_477 = {S_v_3,S_v_2}; // @[RA_Mul.scala 150:21:@739.4]
  assign _T_478 = {_T_477,_T_476}; // @[RA_Mul.scala 150:21:@740.4]
  assign _T_479 = {S_v_5,S_v_4}; // @[RA_Mul.scala 150:21:@741.4]
  assign _T_480 = {S_v_7,S_v_6}; // @[RA_Mul.scala 150:21:@742.4]
  assign _T_481 = {_T_480,_T_479}; // @[RA_Mul.scala 150:21:@743.4]
  assign _T_483 = {SC_v_1,SC_v_0}; // @[RA_Mul.scala 151:23:@746.4]
  assign _T_484 = {SC_v_3,SC_v_2}; // @[RA_Mul.scala 151:23:@747.4]
  assign _T_485 = {_T_484,_T_483}; // @[RA_Mul.scala 151:23:@748.4]
  assign _T_486 = {SC_v_5,SC_v_4}; // @[RA_Mul.scala 151:23:@749.4]
  assign _T_487 = {SC_v_7,SC_v_6}; // @[RA_Mul.scala 151:23:@750.4]
  assign _T_488 = {_T_487,_T_486}; // @[RA_Mul.scala 151:23:@751.4]
  assign io_PP_0 = _T_96 ? 16'h0 : _GEN_3; // @[RA_Mul.scala 126:16:@230.6 RA_Mul.scala 128:16:@235.8 RA_Mul.scala 130:16:@242.10 RA_Mul.scala 132:16:@248.12 RA_Mul.scala 134:16:@256.14 RA_Mul.scala 136:16:@259.14]
  assign io_PP_1 = _T_144 ? 16'h0 : _GEN_10; // @[RA_Mul.scala 126:16:@294.6 RA_Mul.scala 128:16:@299.8 RA_Mul.scala 130:16:@306.10 RA_Mul.scala 132:16:@312.12 RA_Mul.scala 134:16:@320.14 RA_Mul.scala 136:16:@323.14]
  assign io_PP_2 = _T_192 ? 16'h0 : _GEN_17; // @[RA_Mul.scala 126:16:@358.6 RA_Mul.scala 128:16:@363.8 RA_Mul.scala 130:16:@370.10 RA_Mul.scala 132:16:@376.12 RA_Mul.scala 134:16:@384.14 RA_Mul.scala 136:16:@387.14]
  assign io_PP_3 = _T_240 ? 16'h0 : _GEN_24; // @[RA_Mul.scala 126:16:@422.6 RA_Mul.scala 128:16:@427.8 RA_Mul.scala 130:16:@434.10 RA_Mul.scala 132:16:@440.12 RA_Mul.scala 134:16:@448.14 RA_Mul.scala 136:16:@451.14]
  assign io_PP_4 = _T_288 ? 16'h0 : _GEN_31; // @[RA_Mul.scala 126:16:@486.6 RA_Mul.scala 128:16:@491.8 RA_Mul.scala 130:16:@498.10 RA_Mul.scala 132:16:@504.12 RA_Mul.scala 134:16:@512.14 RA_Mul.scala 136:16:@515.14]
  assign io_PP_5 = _T_336 ? 16'h0 : _GEN_38; // @[RA_Mul.scala 126:16:@550.6 RA_Mul.scala 128:16:@555.8 RA_Mul.scala 130:16:@562.10 RA_Mul.scala 132:16:@568.12 RA_Mul.scala 134:16:@576.14 RA_Mul.scala 136:16:@579.14]
  assign io_PP_6 = _T_384 ? 16'h0 : _GEN_45; // @[RA_Mul.scala 126:16:@614.6 RA_Mul.scala 128:16:@619.8 RA_Mul.scala 130:16:@626.10 RA_Mul.scala 132:16:@632.12 RA_Mul.scala 134:16:@640.14 RA_Mul.scala 136:16:@643.14]
  assign io_PP_7 = _T_432 ? 16'h0 : _GEN_52; // @[RA_Mul.scala 126:16:@678.6 RA_Mul.scala 128:16:@683.8 RA_Mul.scala 130:16:@690.10 RA_Mul.scala 132:16:@696.12 RA_Mul.scala 134:16:@704.14 RA_Mul.scala 136:16:@707.14]
  assign io_SC = {_T_488,_T_485}; // @[RA_Mul.scala 151:9:@753.4]
  assign io_S = {_T_481,_T_478}; // @[RA_Mul.scala 150:8:@745.4]
endmodule
module PPLRegs1( // @[:@755.2]
  input         clock, // @[:@756.4]
  input         reset, // @[:@757.4]
  input  [15:0] io_PP_i_0, // @[:@758.4]
  input  [15:0] io_PP_i_1, // @[:@758.4]
  input  [15:0] io_PP_i_2, // @[:@758.4]
  input  [15:0] io_PP_i_3, // @[:@758.4]
  input  [15:0] io_PP_i_4, // @[:@758.4]
  input  [15:0] io_PP_i_5, // @[:@758.4]
  input  [15:0] io_PP_i_6, // @[:@758.4]
  input  [15:0] io_PP_i_7, // @[:@758.4]
  output [15:0] io_PP_o_0, // @[:@758.4]
  output [15:0] io_PP_o_1, // @[:@758.4]
  output [15:0] io_PP_o_2, // @[:@758.4]
  output [15:0] io_PP_o_3, // @[:@758.4]
  output [15:0] io_PP_o_4, // @[:@758.4]
  output [15:0] io_PP_o_5, // @[:@758.4]
  output [15:0] io_PP_o_6, // @[:@758.4]
  output [15:0] io_PP_o_7, // @[:@758.4]
  output [15:0] io_SS_o, // @[:@758.4]
  input  [7:0]  io_SC_i, // @[:@758.4]
  output [7:0]  io_SC_o, // @[:@758.4]
  input  [7:0]  io_S_i, // @[:@758.4]
  output [7:0]  io_S_o // @[:@758.4]
);
  reg [15:0] _T_111_0; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_0;
  reg [15:0] _T_111_1; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_1;
  reg [15:0] _T_111_2; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_2;
  reg [15:0] _T_111_3; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_3;
  reg [15:0] _T_111_4; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_4;
  reg [15:0] _T_111_5; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_5;
  reg [15:0] _T_111_6; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_6;
  reg [15:0] _T_111_7; // @[RA_Mul.scala 671:21:@769.4]
  reg [31:0] _RAND_7;
  reg [15:0] _T_142; // @[RA_Mul.scala 672:21:@786.4]
  reg [31:0] _RAND_8;
  reg [7:0] _T_145; // @[RA_Mul.scala 673:21:@789.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_148; // @[RA_Mul.scala 674:20:@792.4]
  reg [31:0] _RAND_10;
  assign io_PP_o_0 = _T_111_0; // @[RA_Mul.scala 671:11:@778.4]
  assign io_PP_o_1 = _T_111_1; // @[RA_Mul.scala 671:11:@779.4]
  assign io_PP_o_2 = _T_111_2; // @[RA_Mul.scala 671:11:@780.4]
  assign io_PP_o_3 = _T_111_3; // @[RA_Mul.scala 671:11:@781.4]
  assign io_PP_o_4 = _T_111_4; // @[RA_Mul.scala 671:11:@782.4]
  assign io_PP_o_5 = _T_111_5; // @[RA_Mul.scala 671:11:@783.4]
  assign io_PP_o_6 = _T_111_6; // @[RA_Mul.scala 671:11:@784.4]
  assign io_PP_o_7 = _T_111_7; // @[RA_Mul.scala 671:11:@785.4]
  assign io_SS_o = _T_142; // @[RA_Mul.scala 672:11:@788.4]
  assign io_SC_o = _T_145; // @[RA_Mul.scala 673:11:@791.4]
  assign io_S_o = _T_148; // @[RA_Mul.scala 674:10:@794.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_111_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_111_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_111_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_111_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_111_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_111_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_111_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_111_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_142 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_145 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_148 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_111_0 <= 16'h0;
    end else begin
      _T_111_0 <= io_PP_i_0;
    end
    if (reset) begin
      _T_111_1 <= 16'h0;
    end else begin
      _T_111_1 <= io_PP_i_1;
    end
    if (reset) begin
      _T_111_2 <= 16'h0;
    end else begin
      _T_111_2 <= io_PP_i_2;
    end
    if (reset) begin
      _T_111_3 <= 16'h0;
    end else begin
      _T_111_3 <= io_PP_i_3;
    end
    if (reset) begin
      _T_111_4 <= 16'h0;
    end else begin
      _T_111_4 <= io_PP_i_4;
    end
    if (reset) begin
      _T_111_5 <= 16'h0;
    end else begin
      _T_111_5 <= io_PP_i_5;
    end
    if (reset) begin
      _T_111_6 <= 16'h0;
    end else begin
      _T_111_6 <= io_PP_i_6;
    end
    if (reset) begin
      _T_111_7 <= 16'h0;
    end else begin
      _T_111_7 <= io_PP_i_7;
    end
    if (reset) begin
      _T_142 <= 16'h0;
    end else begin
      _T_142 <= 16'haaab;
    end
    if (reset) begin
      _T_145 <= 8'h0;
    end else begin
      _T_145 <= io_SC_i;
    end
    if (reset) begin
      _T_148 <= 8'h0;
    end else begin
      _T_148 <= io_S_i;
    end
  end
endmodule
module HA( // @[:@796.2]
  output  io_s, // @[:@799.4]
  output  io_cout, // @[:@799.4]
  input   io_a, // @[:@799.4]
  input   io_b // @[:@799.4]
);
  assign io_s = io_a ^ io_b; // @[RA_Mul.scala 13:8:@804.4]
  assign io_cout = io_a & io_b; // @[RA_Mul.scala 12:11:@802.4]
endmodule
module FA( // @[:@806.2]
  output  io_s, // @[:@809.4]
  output  io_cout, // @[:@809.4]
  input   io_a, // @[:@809.4]
  input   io_b, // @[:@809.4]
  input   io_cin // @[:@809.4]
);
  wire  _T_15; // @[RA_Mul.scala 36:16:@811.4]
  wire  _T_17; // @[RA_Mul.scala 37:20:@814.4]
  wire  _T_18; // @[RA_Mul.scala 37:36:@815.4]
  wire  _T_19; // @[RA_Mul.scala 37:28:@816.4]
  wire  _T_20; // @[RA_Mul.scala 37:54:@817.4]
  assign _T_15 = io_a ^ io_b; // @[RA_Mul.scala 36:16:@811.4]
  assign _T_17 = io_a & io_b; // @[RA_Mul.scala 37:20:@814.4]
  assign _T_18 = io_a & io_cin; // @[RA_Mul.scala 37:36:@815.4]
  assign _T_19 = _T_17 | _T_18; // @[RA_Mul.scala 37:28:@816.4]
  assign _T_20 = io_b & io_cin; // @[RA_Mul.scala 37:54:@817.4]
  assign io_s = _T_15 ^ io_cin; // @[RA_Mul.scala 36:8:@813.4]
  assign io_cout = _T_19 | _T_20; // @[RA_Mul.scala 37:11:@819.4]
endmodule
module Reduction_1( // @[:@1466.2]
  output        io_matrix_0_0, // @[:@1469.4]
  output        io_matrix_0_1, // @[:@1469.4]
  output        io_matrix_0_2, // @[:@1469.4]
  output        io_matrix_0_3, // @[:@1469.4]
  output        io_matrix_0_4, // @[:@1469.4]
  output        io_matrix_0_5, // @[:@1469.4]
  output        io_matrix_0_6, // @[:@1469.4]
  output        io_matrix_0_7, // @[:@1469.4]
  output        io_matrix_0_8, // @[:@1469.4]
  output        io_matrix_0_9, // @[:@1469.4]
  output        io_matrix_0_10, // @[:@1469.4]
  output        io_matrix_0_11, // @[:@1469.4]
  output        io_matrix_0_12, // @[:@1469.4]
  output        io_matrix_0_13, // @[:@1469.4]
  output        io_matrix_0_14, // @[:@1469.4]
  output        io_matrix_0_15, // @[:@1469.4]
  output        io_matrix_0_16, // @[:@1469.4]
  output        io_matrix_0_17, // @[:@1469.4]
  output        io_matrix_0_18, // @[:@1469.4]
  output        io_matrix_0_19, // @[:@1469.4]
  output        io_matrix_0_20, // @[:@1469.4]
  output        io_matrix_0_21, // @[:@1469.4]
  output        io_matrix_0_22, // @[:@1469.4]
  output        io_matrix_0_23, // @[:@1469.4]
  output        io_matrix_0_24, // @[:@1469.4]
  output        io_matrix_0_25, // @[:@1469.4]
  output        io_matrix_0_26, // @[:@1469.4]
  output        io_matrix_0_27, // @[:@1469.4]
  output        io_matrix_0_28, // @[:@1469.4]
  output        io_matrix_0_29, // @[:@1469.4]
  output        io_matrix_0_30, // @[:@1469.4]
  output        io_matrix_0_31, // @[:@1469.4]
  output        io_matrix_1_1, // @[:@1469.4]
  output        io_matrix_1_3, // @[:@1469.4]
  output        io_matrix_1_4, // @[:@1469.4]
  output        io_matrix_1_5, // @[:@1469.4]
  output        io_matrix_1_6, // @[:@1469.4]
  output        io_matrix_1_7, // @[:@1469.4]
  output        io_matrix_1_8, // @[:@1469.4]
  output        io_matrix_1_9, // @[:@1469.4]
  output        io_matrix_1_10, // @[:@1469.4]
  output        io_matrix_1_11, // @[:@1469.4]
  output        io_matrix_1_12, // @[:@1469.4]
  output        io_matrix_1_13, // @[:@1469.4]
  output        io_matrix_1_14, // @[:@1469.4]
  output        io_matrix_1_15, // @[:@1469.4]
  output        io_matrix_1_16, // @[:@1469.4]
  output        io_matrix_1_17, // @[:@1469.4]
  output        io_matrix_1_18, // @[:@1469.4]
  output        io_matrix_1_19, // @[:@1469.4]
  output        io_matrix_1_20, // @[:@1469.4]
  output        io_matrix_1_21, // @[:@1469.4]
  output        io_matrix_1_22, // @[:@1469.4]
  output        io_matrix_1_23, // @[:@1469.4]
  output        io_matrix_1_24, // @[:@1469.4]
  output        io_matrix_1_25, // @[:@1469.4]
  output        io_matrix_1_26, // @[:@1469.4]
  output        io_matrix_1_27, // @[:@1469.4]
  output        io_matrix_1_28, // @[:@1469.4]
  output        io_matrix_1_29, // @[:@1469.4]
  output        io_matrix_1_30, // @[:@1469.4]
  output        io_matrix_2_3, // @[:@1469.4]
  output        io_matrix_2_6, // @[:@1469.4]
  output        io_matrix_2_7, // @[:@1469.4]
  output        io_matrix_2_8, // @[:@1469.4]
  output        io_matrix_2_9, // @[:@1469.4]
  output        io_matrix_2_10, // @[:@1469.4]
  output        io_matrix_2_11, // @[:@1469.4]
  output        io_matrix_2_12, // @[:@1469.4]
  output        io_matrix_2_13, // @[:@1469.4]
  output        io_matrix_2_14, // @[:@1469.4]
  output        io_matrix_2_15, // @[:@1469.4]
  output        io_matrix_2_16, // @[:@1469.4]
  output        io_matrix_2_17, // @[:@1469.4]
  output        io_matrix_2_18, // @[:@1469.4]
  output        io_matrix_2_19, // @[:@1469.4]
  output        io_matrix_2_20, // @[:@1469.4]
  output        io_matrix_2_21, // @[:@1469.4]
  output        io_matrix_2_22, // @[:@1469.4]
  output        io_matrix_2_23, // @[:@1469.4]
  output        io_matrix_2_24, // @[:@1469.4]
  output        io_matrix_2_25, // @[:@1469.4]
  output        io_matrix_2_26, // @[:@1469.4]
  output        io_matrix_2_29, // @[:@1469.4]
  output        io_matrix_3_6, // @[:@1469.4]
  output        io_matrix_3_9, // @[:@1469.4]
  output        io_matrix_3_10, // @[:@1469.4]
  output        io_matrix_3_11, // @[:@1469.4]
  output        io_matrix_3_12, // @[:@1469.4]
  output        io_matrix_3_13, // @[:@1469.4]
  output        io_matrix_3_14, // @[:@1469.4]
  output        io_matrix_3_15, // @[:@1469.4]
  output        io_matrix_3_16, // @[:@1469.4]
  output        io_matrix_3_17, // @[:@1469.4]
  output        io_matrix_3_18, // @[:@1469.4]
  output        io_matrix_3_19, // @[:@1469.4]
  output        io_matrix_3_20, // @[:@1469.4]
  output        io_matrix_3_21, // @[:@1469.4]
  output        io_matrix_3_22, // @[:@1469.4]
  output        io_matrix_3_23, // @[:@1469.4]
  output        io_matrix_3_24, // @[:@1469.4]
  output        io_matrix_4_9, // @[:@1469.4]
  output        io_matrix_4_12, // @[:@1469.4]
  output        io_matrix_4_13, // @[:@1469.4]
  output        io_matrix_4_14, // @[:@1469.4]
  output        io_matrix_4_15, // @[:@1469.4]
  output        io_matrix_4_16, // @[:@1469.4]
  output        io_matrix_4_17, // @[:@1469.4]
  output        io_matrix_4_18, // @[:@1469.4]
  output        io_matrix_4_19, // @[:@1469.4]
  output        io_matrix_4_20, // @[:@1469.4]
  output        io_matrix_4_23, // @[:@1469.4]
  output        io_matrix_5_12, // @[:@1469.4]
  output        io_matrix_5_15, // @[:@1469.4]
  output        io_matrix_5_16, // @[:@1469.4]
  output        io_matrix_5_17, // @[:@1469.4]
  output        io_matrix_5_18, // @[:@1469.4]
  output        io_matrix_5_19, // @[:@1469.4]
  input  [15:0] io_PP_0, // @[:@1469.4]
  input  [15:0] io_PP_1, // @[:@1469.4]
  input  [15:0] io_PP_2, // @[:@1469.4]
  input  [15:0] io_PP_3, // @[:@1469.4]
  input  [15:0] io_PP_4, // @[:@1469.4]
  input  [15:0] io_PP_5, // @[:@1469.4]
  input  [15:0] io_PP_6, // @[:@1469.4]
  input  [15:0] io_PP_7, // @[:@1469.4]
  input  [15:0] io_SS, // @[:@1469.4]
  input  [7:0]  io_SC, // @[:@1469.4]
  input  [7:0]  io_S // @[:@1469.4]
);
  wire  HA_io_s; // @[RA_Mul.scala 19:21:@1473.4]
  wire  HA_io_cout; // @[RA_Mul.scala 19:21:@1473.4]
  wire  HA_io_a; // @[RA_Mul.scala 19:21:@1473.4]
  wire  HA_io_b; // @[RA_Mul.scala 19:21:@1473.4]
  wire  FA_io_s; // @[RA_Mul.scala 43:21:@1494.4]
  wire  FA_io_cout; // @[RA_Mul.scala 43:21:@1494.4]
  wire  FA_io_a; // @[RA_Mul.scala 43:21:@1494.4]
  wire  FA_io_b; // @[RA_Mul.scala 43:21:@1494.4]
  wire  FA_io_cin; // @[RA_Mul.scala 43:21:@1494.4]
  wire  FA_1_io_s; // @[RA_Mul.scala 43:21:@1517.4]
  wire  FA_1_io_cout; // @[RA_Mul.scala 43:21:@1517.4]
  wire  FA_1_io_a; // @[RA_Mul.scala 43:21:@1517.4]
  wire  FA_1_io_b; // @[RA_Mul.scala 43:21:@1517.4]
  wire  FA_1_io_cin; // @[RA_Mul.scala 43:21:@1517.4]
  wire  FA_2_io_s; // @[RA_Mul.scala 43:21:@1534.4]
  wire  FA_2_io_cout; // @[RA_Mul.scala 43:21:@1534.4]
  wire  FA_2_io_a; // @[RA_Mul.scala 43:21:@1534.4]
  wire  FA_2_io_b; // @[RA_Mul.scala 43:21:@1534.4]
  wire  FA_2_io_cin; // @[RA_Mul.scala 43:21:@1534.4]
  wire  FA_3_io_s; // @[RA_Mul.scala 43:21:@1549.4]
  wire  FA_3_io_cout; // @[RA_Mul.scala 43:21:@1549.4]
  wire  FA_3_io_a; // @[RA_Mul.scala 43:21:@1549.4]
  wire  FA_3_io_b; // @[RA_Mul.scala 43:21:@1549.4]
  wire  FA_3_io_cin; // @[RA_Mul.scala 43:21:@1549.4]
  wire  FA_4_io_s; // @[RA_Mul.scala 43:21:@1566.4]
  wire  FA_4_io_cout; // @[RA_Mul.scala 43:21:@1566.4]
  wire  FA_4_io_a; // @[RA_Mul.scala 43:21:@1566.4]
  wire  FA_4_io_b; // @[RA_Mul.scala 43:21:@1566.4]
  wire  FA_4_io_cin; // @[RA_Mul.scala 43:21:@1566.4]
  wire  FA_5_io_s; // @[RA_Mul.scala 43:21:@1582.4]
  wire  FA_5_io_cout; // @[RA_Mul.scala 43:21:@1582.4]
  wire  FA_5_io_a; // @[RA_Mul.scala 43:21:@1582.4]
  wire  FA_5_io_b; // @[RA_Mul.scala 43:21:@1582.4]
  wire  FA_5_io_cin; // @[RA_Mul.scala 43:21:@1582.4]
  wire  FA_6_io_s; // @[RA_Mul.scala 43:21:@1593.4]
  wire  FA_6_io_cout; // @[RA_Mul.scala 43:21:@1593.4]
  wire  FA_6_io_a; // @[RA_Mul.scala 43:21:@1593.4]
  wire  FA_6_io_b; // @[RA_Mul.scala 43:21:@1593.4]
  wire  FA_6_io_cin; // @[RA_Mul.scala 43:21:@1593.4]
  wire  FA_7_io_s; // @[RA_Mul.scala 43:21:@1607.4]
  wire  FA_7_io_cout; // @[RA_Mul.scala 43:21:@1607.4]
  wire  FA_7_io_a; // @[RA_Mul.scala 43:21:@1607.4]
  wire  FA_7_io_b; // @[RA_Mul.scala 43:21:@1607.4]
  wire  FA_7_io_cin; // @[RA_Mul.scala 43:21:@1607.4]
  wire  FA_8_io_s; // @[RA_Mul.scala 43:21:@1623.4]
  wire  FA_8_io_cout; // @[RA_Mul.scala 43:21:@1623.4]
  wire  FA_8_io_a; // @[RA_Mul.scala 43:21:@1623.4]
  wire  FA_8_io_b; // @[RA_Mul.scala 43:21:@1623.4]
  wire  FA_8_io_cin; // @[RA_Mul.scala 43:21:@1623.4]
  wire  FA_9_io_s; // @[RA_Mul.scala 43:21:@1634.4]
  wire  FA_9_io_cout; // @[RA_Mul.scala 43:21:@1634.4]
  wire  FA_9_io_a; // @[RA_Mul.scala 43:21:@1634.4]
  wire  FA_9_io_b; // @[RA_Mul.scala 43:21:@1634.4]
  wire  FA_9_io_cin; // @[RA_Mul.scala 43:21:@1634.4]
  wire  FA_10_io_s; // @[RA_Mul.scala 43:21:@1649.4]
  wire  FA_10_io_cout; // @[RA_Mul.scala 43:21:@1649.4]
  wire  FA_10_io_a; // @[RA_Mul.scala 43:21:@1649.4]
  wire  FA_10_io_b; // @[RA_Mul.scala 43:21:@1649.4]
  wire  FA_10_io_cin; // @[RA_Mul.scala 43:21:@1649.4]
  wire  FA_11_io_s; // @[RA_Mul.scala 43:21:@1660.4]
  wire  FA_11_io_cout; // @[RA_Mul.scala 43:21:@1660.4]
  wire  FA_11_io_a; // @[RA_Mul.scala 43:21:@1660.4]
  wire  FA_11_io_b; // @[RA_Mul.scala 43:21:@1660.4]
  wire  FA_11_io_cin; // @[RA_Mul.scala 43:21:@1660.4]
  wire  FA_12_io_s; // @[RA_Mul.scala 43:21:@1673.4]
  wire  FA_12_io_cout; // @[RA_Mul.scala 43:21:@1673.4]
  wire  FA_12_io_a; // @[RA_Mul.scala 43:21:@1673.4]
  wire  FA_12_io_b; // @[RA_Mul.scala 43:21:@1673.4]
  wire  FA_12_io_cin; // @[RA_Mul.scala 43:21:@1673.4]
  wire  FA_13_io_s; // @[RA_Mul.scala 43:21:@1684.4]
  wire  FA_13_io_cout; // @[RA_Mul.scala 43:21:@1684.4]
  wire  FA_13_io_a; // @[RA_Mul.scala 43:21:@1684.4]
  wire  FA_13_io_b; // @[RA_Mul.scala 43:21:@1684.4]
  wire  FA_13_io_cin; // @[RA_Mul.scala 43:21:@1684.4]
  wire  FA_14_io_s; // @[RA_Mul.scala 43:21:@1699.4]
  wire  FA_14_io_cout; // @[RA_Mul.scala 43:21:@1699.4]
  wire  FA_14_io_a; // @[RA_Mul.scala 43:21:@1699.4]
  wire  FA_14_io_b; // @[RA_Mul.scala 43:21:@1699.4]
  wire  FA_14_io_cin; // @[RA_Mul.scala 43:21:@1699.4]
  wire  FA_15_io_s; // @[RA_Mul.scala 43:21:@1710.4]
  wire  FA_15_io_cout; // @[RA_Mul.scala 43:21:@1710.4]
  wire  FA_15_io_a; // @[RA_Mul.scala 43:21:@1710.4]
  wire  FA_15_io_b; // @[RA_Mul.scala 43:21:@1710.4]
  wire  FA_15_io_cin; // @[RA_Mul.scala 43:21:@1710.4]
  wire  FA_16_io_s; // @[RA_Mul.scala 43:21:@1724.4]
  wire  FA_16_io_cout; // @[RA_Mul.scala 43:21:@1724.4]
  wire  FA_16_io_a; // @[RA_Mul.scala 43:21:@1724.4]
  wire  FA_16_io_b; // @[RA_Mul.scala 43:21:@1724.4]
  wire  FA_16_io_cin; // @[RA_Mul.scala 43:21:@1724.4]
  wire  FA_17_io_s; // @[RA_Mul.scala 43:21:@1735.4]
  wire  FA_17_io_cout; // @[RA_Mul.scala 43:21:@1735.4]
  wire  FA_17_io_a; // @[RA_Mul.scala 43:21:@1735.4]
  wire  FA_17_io_b; // @[RA_Mul.scala 43:21:@1735.4]
  wire  FA_17_io_cin; // @[RA_Mul.scala 43:21:@1735.4]
  wire  FA_18_io_s; // @[RA_Mul.scala 43:21:@1746.4]
  wire  FA_18_io_cout; // @[RA_Mul.scala 43:21:@1746.4]
  wire  FA_18_io_a; // @[RA_Mul.scala 43:21:@1746.4]
  wire  FA_18_io_b; // @[RA_Mul.scala 43:21:@1746.4]
  wire  FA_18_io_cin; // @[RA_Mul.scala 43:21:@1746.4]
  wire  FA_19_io_s; // @[RA_Mul.scala 43:21:@1758.4]
  wire  FA_19_io_cout; // @[RA_Mul.scala 43:21:@1758.4]
  wire  FA_19_io_a; // @[RA_Mul.scala 43:21:@1758.4]
  wire  FA_19_io_b; // @[RA_Mul.scala 43:21:@1758.4]
  wire  FA_19_io_cin; // @[RA_Mul.scala 43:21:@1758.4]
  wire  FA_20_io_s; // @[RA_Mul.scala 43:21:@1769.4]
  wire  FA_20_io_cout; // @[RA_Mul.scala 43:21:@1769.4]
  wire  FA_20_io_a; // @[RA_Mul.scala 43:21:@1769.4]
  wire  FA_20_io_b; // @[RA_Mul.scala 43:21:@1769.4]
  wire  FA_20_io_cin; // @[RA_Mul.scala 43:21:@1769.4]
  wire  HA_1_io_s; // @[RA_Mul.scala 19:21:@1779.4]
  wire  HA_1_io_cout; // @[RA_Mul.scala 19:21:@1779.4]
  wire  HA_1_io_a; // @[RA_Mul.scala 19:21:@1779.4]
  wire  HA_1_io_b; // @[RA_Mul.scala 19:21:@1779.4]
  wire  FA_21_io_s; // @[RA_Mul.scala 43:21:@1789.4]
  wire  FA_21_io_cout; // @[RA_Mul.scala 43:21:@1789.4]
  wire  FA_21_io_a; // @[RA_Mul.scala 43:21:@1789.4]
  wire  FA_21_io_b; // @[RA_Mul.scala 43:21:@1789.4]
  wire  FA_21_io_cin; // @[RA_Mul.scala 43:21:@1789.4]
  wire  FA_22_io_s; // @[RA_Mul.scala 43:21:@1800.4]
  wire  FA_22_io_cout; // @[RA_Mul.scala 43:21:@1800.4]
  wire  FA_22_io_a; // @[RA_Mul.scala 43:21:@1800.4]
  wire  FA_22_io_b; // @[RA_Mul.scala 43:21:@1800.4]
  wire  FA_22_io_cin; // @[RA_Mul.scala 43:21:@1800.4]
  wire  FA_23_io_s; // @[RA_Mul.scala 43:21:@1811.4]
  wire  FA_23_io_cout; // @[RA_Mul.scala 43:21:@1811.4]
  wire  FA_23_io_a; // @[RA_Mul.scala 43:21:@1811.4]
  wire  FA_23_io_b; // @[RA_Mul.scala 43:21:@1811.4]
  wire  FA_23_io_cin; // @[RA_Mul.scala 43:21:@1811.4]
  wire  FA_24_io_s; // @[RA_Mul.scala 43:21:@1822.4]
  wire  FA_24_io_cout; // @[RA_Mul.scala 43:21:@1822.4]
  wire  FA_24_io_a; // @[RA_Mul.scala 43:21:@1822.4]
  wire  FA_24_io_b; // @[RA_Mul.scala 43:21:@1822.4]
  wire  FA_24_io_cin; // @[RA_Mul.scala 43:21:@1822.4]
  wire  FA_25_io_s; // @[RA_Mul.scala 43:21:@1833.4]
  wire  FA_25_io_cout; // @[RA_Mul.scala 43:21:@1833.4]
  wire  FA_25_io_a; // @[RA_Mul.scala 43:21:@1833.4]
  wire  FA_25_io_b; // @[RA_Mul.scala 43:21:@1833.4]
  wire  FA_25_io_cin; // @[RA_Mul.scala 43:21:@1833.4]
  wire  HA_2_io_s; // @[RA_Mul.scala 19:21:@1843.4]
  wire  HA_2_io_cout; // @[RA_Mul.scala 19:21:@1843.4]
  wire  HA_2_io_a; // @[RA_Mul.scala 19:21:@1843.4]
  wire  HA_2_io_b; // @[RA_Mul.scala 19:21:@1843.4]
  wire  FA_26_io_s; // @[RA_Mul.scala 43:21:@1853.4]
  wire  FA_26_io_cout; // @[RA_Mul.scala 43:21:@1853.4]
  wire  FA_26_io_a; // @[RA_Mul.scala 43:21:@1853.4]
  wire  FA_26_io_b; // @[RA_Mul.scala 43:21:@1853.4]
  wire  FA_26_io_cin; // @[RA_Mul.scala 43:21:@1853.4]
  wire  FA_27_io_s; // @[RA_Mul.scala 43:21:@1864.4]
  wire  FA_27_io_cout; // @[RA_Mul.scala 43:21:@1864.4]
  wire  FA_27_io_a; // @[RA_Mul.scala 43:21:@1864.4]
  wire  FA_27_io_b; // @[RA_Mul.scala 43:21:@1864.4]
  wire  FA_27_io_cin; // @[RA_Mul.scala 43:21:@1864.4]
  wire  HA_3_io_s; // @[RA_Mul.scala 19:21:@1874.4]
  wire  HA_3_io_cout; // @[RA_Mul.scala 19:21:@1874.4]
  wire  HA_3_io_a; // @[RA_Mul.scala 19:21:@1874.4]
  wire  HA_3_io_b; // @[RA_Mul.scala 19:21:@1874.4]
  wire  FA_28_io_s; // @[RA_Mul.scala 43:21:@1884.4]
  wire  FA_28_io_cout; // @[RA_Mul.scala 43:21:@1884.4]
  wire  FA_28_io_a; // @[RA_Mul.scala 43:21:@1884.4]
  wire  FA_28_io_b; // @[RA_Mul.scala 43:21:@1884.4]
  wire  FA_28_io_cin; // @[RA_Mul.scala 43:21:@1884.4]
  wire  FA_29_io_s; // @[RA_Mul.scala 43:21:@1895.4]
  wire  FA_29_io_cout; // @[RA_Mul.scala 43:21:@1895.4]
  wire  FA_29_io_a; // @[RA_Mul.scala 43:21:@1895.4]
  wire  FA_29_io_b; // @[RA_Mul.scala 43:21:@1895.4]
  wire  FA_29_io_cin; // @[RA_Mul.scala 43:21:@1895.4]
  wire  FA_30_io_s; // @[RA_Mul.scala 43:21:@1908.4]
  wire  FA_30_io_cout; // @[RA_Mul.scala 43:21:@1908.4]
  wire  FA_30_io_a; // @[RA_Mul.scala 43:21:@1908.4]
  wire  FA_30_io_b; // @[RA_Mul.scala 43:21:@1908.4]
  wire  FA_30_io_cin; // @[RA_Mul.scala 43:21:@1908.4]
  wire  FA_31_io_s; // @[RA_Mul.scala 43:21:@1919.4]
  wire  FA_31_io_cout; // @[RA_Mul.scala 43:21:@1919.4]
  wire  FA_31_io_a; // @[RA_Mul.scala 43:21:@1919.4]
  wire  FA_31_io_b; // @[RA_Mul.scala 43:21:@1919.4]
  wire  FA_31_io_cin; // @[RA_Mul.scala 43:21:@1919.4]
  wire  FA_32_io_s; // @[RA_Mul.scala 43:21:@1933.4]
  wire  FA_32_io_cout; // @[RA_Mul.scala 43:21:@1933.4]
  wire  FA_32_io_a; // @[RA_Mul.scala 43:21:@1933.4]
  wire  FA_32_io_b; // @[RA_Mul.scala 43:21:@1933.4]
  wire  FA_32_io_cin; // @[RA_Mul.scala 43:21:@1933.4]
  wire  FA_33_io_s; // @[RA_Mul.scala 43:21:@1944.4]
  wire  FA_33_io_cout; // @[RA_Mul.scala 43:21:@1944.4]
  wire  FA_33_io_a; // @[RA_Mul.scala 43:21:@1944.4]
  wire  FA_33_io_b; // @[RA_Mul.scala 43:21:@1944.4]
  wire  FA_33_io_cin; // @[RA_Mul.scala 43:21:@1944.4]
  wire  FA_34_io_s; // @[RA_Mul.scala 43:21:@1957.4]
  wire  FA_34_io_cout; // @[RA_Mul.scala 43:21:@1957.4]
  wire  FA_34_io_a; // @[RA_Mul.scala 43:21:@1957.4]
  wire  FA_34_io_b; // @[RA_Mul.scala 43:21:@1957.4]
  wire  FA_34_io_cin; // @[RA_Mul.scala 43:21:@1957.4]
  wire  FA_35_io_s; // @[RA_Mul.scala 43:21:@1968.4]
  wire  FA_35_io_cout; // @[RA_Mul.scala 43:21:@1968.4]
  wire  FA_35_io_a; // @[RA_Mul.scala 43:21:@1968.4]
  wire  FA_35_io_b; // @[RA_Mul.scala 43:21:@1968.4]
  wire  FA_35_io_cin; // @[RA_Mul.scala 43:21:@1968.4]
  wire  FA_36_io_s; // @[RA_Mul.scala 43:21:@1981.4]
  wire  FA_36_io_cout; // @[RA_Mul.scala 43:21:@1981.4]
  wire  FA_36_io_a; // @[RA_Mul.scala 43:21:@1981.4]
  wire  FA_36_io_b; // @[RA_Mul.scala 43:21:@1981.4]
  wire  FA_36_io_cin; // @[RA_Mul.scala 43:21:@1981.4]
  wire  FA_37_io_s; // @[RA_Mul.scala 43:21:@1997.4]
  wire  FA_37_io_cout; // @[RA_Mul.scala 43:21:@1997.4]
  wire  FA_37_io_a; // @[RA_Mul.scala 43:21:@1997.4]
  wire  FA_37_io_b; // @[RA_Mul.scala 43:21:@1997.4]
  wire  FA_37_io_cin; // @[RA_Mul.scala 43:21:@1997.4]
  wire  FA_38_io_s; // @[RA_Mul.scala 43:21:@2014.4]
  wire  FA_38_io_cout; // @[RA_Mul.scala 43:21:@2014.4]
  wire  FA_38_io_a; // @[RA_Mul.scala 43:21:@2014.4]
  wire  FA_38_io_b; // @[RA_Mul.scala 43:21:@2014.4]
  wire  FA_38_io_cin; // @[RA_Mul.scala 43:21:@2014.4]
  wire  FA_39_io_s; // @[RA_Mul.scala 43:21:@2030.4]
  wire  FA_39_io_cout; // @[RA_Mul.scala 43:21:@2030.4]
  wire  FA_39_io_a; // @[RA_Mul.scala 43:21:@2030.4]
  wire  FA_39_io_b; // @[RA_Mul.scala 43:21:@2030.4]
  wire  FA_39_io_cin; // @[RA_Mul.scala 43:21:@2030.4]
  wire  FA_40_io_s; // @[RA_Mul.scala 43:21:@2046.4]
  wire  FA_40_io_cout; // @[RA_Mul.scala 43:21:@2046.4]
  wire  FA_40_io_a; // @[RA_Mul.scala 43:21:@2046.4]
  wire  FA_40_io_b; // @[RA_Mul.scala 43:21:@2046.4]
  wire  FA_40_io_cin; // @[RA_Mul.scala 43:21:@2046.4]
  wire  FA_41_io_s; // @[RA_Mul.scala 43:21:@2061.4]
  wire  FA_41_io_cout; // @[RA_Mul.scala 43:21:@2061.4]
  wire  FA_41_io_a; // @[RA_Mul.scala 43:21:@2061.4]
  wire  FA_41_io_b; // @[RA_Mul.scala 43:21:@2061.4]
  wire  FA_41_io_cin; // @[RA_Mul.scala 43:21:@2061.4]
  HA HA ( // @[RA_Mul.scala 19:21:@1473.4]
    .io_s(HA_io_s),
    .io_cout(HA_io_cout),
    .io_a(HA_io_a),
    .io_b(HA_io_b)
  );
  FA FA ( // @[RA_Mul.scala 43:21:@1494.4]
    .io_s(FA_io_s),
    .io_cout(FA_io_cout),
    .io_a(FA_io_a),
    .io_b(FA_io_b),
    .io_cin(FA_io_cin)
  );
  FA FA_1 ( // @[RA_Mul.scala 43:21:@1517.4]
    .io_s(FA_1_io_s),
    .io_cout(FA_1_io_cout),
    .io_a(FA_1_io_a),
    .io_b(FA_1_io_b),
    .io_cin(FA_1_io_cin)
  );
  FA FA_2 ( // @[RA_Mul.scala 43:21:@1534.4]
    .io_s(FA_2_io_s),
    .io_cout(FA_2_io_cout),
    .io_a(FA_2_io_a),
    .io_b(FA_2_io_b),
    .io_cin(FA_2_io_cin)
  );
  FA FA_3 ( // @[RA_Mul.scala 43:21:@1549.4]
    .io_s(FA_3_io_s),
    .io_cout(FA_3_io_cout),
    .io_a(FA_3_io_a),
    .io_b(FA_3_io_b),
    .io_cin(FA_3_io_cin)
  );
  FA FA_4 ( // @[RA_Mul.scala 43:21:@1566.4]
    .io_s(FA_4_io_s),
    .io_cout(FA_4_io_cout),
    .io_a(FA_4_io_a),
    .io_b(FA_4_io_b),
    .io_cin(FA_4_io_cin)
  );
  FA FA_5 ( // @[RA_Mul.scala 43:21:@1582.4]
    .io_s(FA_5_io_s),
    .io_cout(FA_5_io_cout),
    .io_a(FA_5_io_a),
    .io_b(FA_5_io_b),
    .io_cin(FA_5_io_cin)
  );
  FA FA_6 ( // @[RA_Mul.scala 43:21:@1593.4]
    .io_s(FA_6_io_s),
    .io_cout(FA_6_io_cout),
    .io_a(FA_6_io_a),
    .io_b(FA_6_io_b),
    .io_cin(FA_6_io_cin)
  );
  FA FA_7 ( // @[RA_Mul.scala 43:21:@1607.4]
    .io_s(FA_7_io_s),
    .io_cout(FA_7_io_cout),
    .io_a(FA_7_io_a),
    .io_b(FA_7_io_b),
    .io_cin(FA_7_io_cin)
  );
  FA FA_8 ( // @[RA_Mul.scala 43:21:@1623.4]
    .io_s(FA_8_io_s),
    .io_cout(FA_8_io_cout),
    .io_a(FA_8_io_a),
    .io_b(FA_8_io_b),
    .io_cin(FA_8_io_cin)
  );
  FA FA_9 ( // @[RA_Mul.scala 43:21:@1634.4]
    .io_s(FA_9_io_s),
    .io_cout(FA_9_io_cout),
    .io_a(FA_9_io_a),
    .io_b(FA_9_io_b),
    .io_cin(FA_9_io_cin)
  );
  FA FA_10 ( // @[RA_Mul.scala 43:21:@1649.4]
    .io_s(FA_10_io_s),
    .io_cout(FA_10_io_cout),
    .io_a(FA_10_io_a),
    .io_b(FA_10_io_b),
    .io_cin(FA_10_io_cin)
  );
  FA FA_11 ( // @[RA_Mul.scala 43:21:@1660.4]
    .io_s(FA_11_io_s),
    .io_cout(FA_11_io_cout),
    .io_a(FA_11_io_a),
    .io_b(FA_11_io_b),
    .io_cin(FA_11_io_cin)
  );
  FA FA_12 ( // @[RA_Mul.scala 43:21:@1673.4]
    .io_s(FA_12_io_s),
    .io_cout(FA_12_io_cout),
    .io_a(FA_12_io_a),
    .io_b(FA_12_io_b),
    .io_cin(FA_12_io_cin)
  );
  FA FA_13 ( // @[RA_Mul.scala 43:21:@1684.4]
    .io_s(FA_13_io_s),
    .io_cout(FA_13_io_cout),
    .io_a(FA_13_io_a),
    .io_b(FA_13_io_b),
    .io_cin(FA_13_io_cin)
  );
  FA FA_14 ( // @[RA_Mul.scala 43:21:@1699.4]
    .io_s(FA_14_io_s),
    .io_cout(FA_14_io_cout),
    .io_a(FA_14_io_a),
    .io_b(FA_14_io_b),
    .io_cin(FA_14_io_cin)
  );
  FA FA_15 ( // @[RA_Mul.scala 43:21:@1710.4]
    .io_s(FA_15_io_s),
    .io_cout(FA_15_io_cout),
    .io_a(FA_15_io_a),
    .io_b(FA_15_io_b),
    .io_cin(FA_15_io_cin)
  );
  FA FA_16 ( // @[RA_Mul.scala 43:21:@1724.4]
    .io_s(FA_16_io_s),
    .io_cout(FA_16_io_cout),
    .io_a(FA_16_io_a),
    .io_b(FA_16_io_b),
    .io_cin(FA_16_io_cin)
  );
  FA FA_17 ( // @[RA_Mul.scala 43:21:@1735.4]
    .io_s(FA_17_io_s),
    .io_cout(FA_17_io_cout),
    .io_a(FA_17_io_a),
    .io_b(FA_17_io_b),
    .io_cin(FA_17_io_cin)
  );
  FA FA_18 ( // @[RA_Mul.scala 43:21:@1746.4]
    .io_s(FA_18_io_s),
    .io_cout(FA_18_io_cout),
    .io_a(FA_18_io_a),
    .io_b(FA_18_io_b),
    .io_cin(FA_18_io_cin)
  );
  FA FA_19 ( // @[RA_Mul.scala 43:21:@1758.4]
    .io_s(FA_19_io_s),
    .io_cout(FA_19_io_cout),
    .io_a(FA_19_io_a),
    .io_b(FA_19_io_b),
    .io_cin(FA_19_io_cin)
  );
  FA FA_20 ( // @[RA_Mul.scala 43:21:@1769.4]
    .io_s(FA_20_io_s),
    .io_cout(FA_20_io_cout),
    .io_a(FA_20_io_a),
    .io_b(FA_20_io_b),
    .io_cin(FA_20_io_cin)
  );
  HA HA_1 ( // @[RA_Mul.scala 19:21:@1779.4]
    .io_s(HA_1_io_s),
    .io_cout(HA_1_io_cout),
    .io_a(HA_1_io_a),
    .io_b(HA_1_io_b)
  );
  FA FA_21 ( // @[RA_Mul.scala 43:21:@1789.4]
    .io_s(FA_21_io_s),
    .io_cout(FA_21_io_cout),
    .io_a(FA_21_io_a),
    .io_b(FA_21_io_b),
    .io_cin(FA_21_io_cin)
  );
  FA FA_22 ( // @[RA_Mul.scala 43:21:@1800.4]
    .io_s(FA_22_io_s),
    .io_cout(FA_22_io_cout),
    .io_a(FA_22_io_a),
    .io_b(FA_22_io_b),
    .io_cin(FA_22_io_cin)
  );
  FA FA_23 ( // @[RA_Mul.scala 43:21:@1811.4]
    .io_s(FA_23_io_s),
    .io_cout(FA_23_io_cout),
    .io_a(FA_23_io_a),
    .io_b(FA_23_io_b),
    .io_cin(FA_23_io_cin)
  );
  FA FA_24 ( // @[RA_Mul.scala 43:21:@1822.4]
    .io_s(FA_24_io_s),
    .io_cout(FA_24_io_cout),
    .io_a(FA_24_io_a),
    .io_b(FA_24_io_b),
    .io_cin(FA_24_io_cin)
  );
  FA FA_25 ( // @[RA_Mul.scala 43:21:@1833.4]
    .io_s(FA_25_io_s),
    .io_cout(FA_25_io_cout),
    .io_a(FA_25_io_a),
    .io_b(FA_25_io_b),
    .io_cin(FA_25_io_cin)
  );
  HA HA_2 ( // @[RA_Mul.scala 19:21:@1843.4]
    .io_s(HA_2_io_s),
    .io_cout(HA_2_io_cout),
    .io_a(HA_2_io_a),
    .io_b(HA_2_io_b)
  );
  FA FA_26 ( // @[RA_Mul.scala 43:21:@1853.4]
    .io_s(FA_26_io_s),
    .io_cout(FA_26_io_cout),
    .io_a(FA_26_io_a),
    .io_b(FA_26_io_b),
    .io_cin(FA_26_io_cin)
  );
  FA FA_27 ( // @[RA_Mul.scala 43:21:@1864.4]
    .io_s(FA_27_io_s),
    .io_cout(FA_27_io_cout),
    .io_a(FA_27_io_a),
    .io_b(FA_27_io_b),
    .io_cin(FA_27_io_cin)
  );
  HA HA_3 ( // @[RA_Mul.scala 19:21:@1874.4]
    .io_s(HA_3_io_s),
    .io_cout(HA_3_io_cout),
    .io_a(HA_3_io_a),
    .io_b(HA_3_io_b)
  );
  FA FA_28 ( // @[RA_Mul.scala 43:21:@1884.4]
    .io_s(FA_28_io_s),
    .io_cout(FA_28_io_cout),
    .io_a(FA_28_io_a),
    .io_b(FA_28_io_b),
    .io_cin(FA_28_io_cin)
  );
  FA FA_29 ( // @[RA_Mul.scala 43:21:@1895.4]
    .io_s(FA_29_io_s),
    .io_cout(FA_29_io_cout),
    .io_a(FA_29_io_a),
    .io_b(FA_29_io_b),
    .io_cin(FA_29_io_cin)
  );
  FA FA_30 ( // @[RA_Mul.scala 43:21:@1908.4]
    .io_s(FA_30_io_s),
    .io_cout(FA_30_io_cout),
    .io_a(FA_30_io_a),
    .io_b(FA_30_io_b),
    .io_cin(FA_30_io_cin)
  );
  FA FA_31 ( // @[RA_Mul.scala 43:21:@1919.4]
    .io_s(FA_31_io_s),
    .io_cout(FA_31_io_cout),
    .io_a(FA_31_io_a),
    .io_b(FA_31_io_b),
    .io_cin(FA_31_io_cin)
  );
  FA FA_32 ( // @[RA_Mul.scala 43:21:@1933.4]
    .io_s(FA_32_io_s),
    .io_cout(FA_32_io_cout),
    .io_a(FA_32_io_a),
    .io_b(FA_32_io_b),
    .io_cin(FA_32_io_cin)
  );
  FA FA_33 ( // @[RA_Mul.scala 43:21:@1944.4]
    .io_s(FA_33_io_s),
    .io_cout(FA_33_io_cout),
    .io_a(FA_33_io_a),
    .io_b(FA_33_io_b),
    .io_cin(FA_33_io_cin)
  );
  FA FA_34 ( // @[RA_Mul.scala 43:21:@1957.4]
    .io_s(FA_34_io_s),
    .io_cout(FA_34_io_cout),
    .io_a(FA_34_io_a),
    .io_b(FA_34_io_b),
    .io_cin(FA_34_io_cin)
  );
  FA FA_35 ( // @[RA_Mul.scala 43:21:@1968.4]
    .io_s(FA_35_io_s),
    .io_cout(FA_35_io_cout),
    .io_a(FA_35_io_a),
    .io_b(FA_35_io_b),
    .io_cin(FA_35_io_cin)
  );
  FA FA_36 ( // @[RA_Mul.scala 43:21:@1981.4]
    .io_s(FA_36_io_s),
    .io_cout(FA_36_io_cout),
    .io_a(FA_36_io_a),
    .io_b(FA_36_io_b),
    .io_cin(FA_36_io_cin)
  );
  FA FA_37 ( // @[RA_Mul.scala 43:21:@1997.4]
    .io_s(FA_37_io_s),
    .io_cout(FA_37_io_cout),
    .io_a(FA_37_io_a),
    .io_b(FA_37_io_b),
    .io_cin(FA_37_io_cin)
  );
  FA FA_38 ( // @[RA_Mul.scala 43:21:@2014.4]
    .io_s(FA_38_io_s),
    .io_cout(FA_38_io_cout),
    .io_a(FA_38_io_a),
    .io_b(FA_38_io_b),
    .io_cin(FA_38_io_cin)
  );
  FA FA_39 ( // @[RA_Mul.scala 43:21:@2030.4]
    .io_s(FA_39_io_s),
    .io_cout(FA_39_io_cout),
    .io_a(FA_39_io_a),
    .io_b(FA_39_io_b),
    .io_cin(FA_39_io_cin)
  );
  FA FA_40 ( // @[RA_Mul.scala 43:21:@2046.4]
    .io_s(FA_40_io_s),
    .io_cout(FA_40_io_cout),
    .io_a(FA_40_io_a),
    .io_b(FA_40_io_b),
    .io_cin(FA_40_io_cin)
  );
  FA FA_41 ( // @[RA_Mul.scala 43:21:@2061.4]
    .io_s(FA_41_io_s),
    .io_cout(FA_41_io_cout),
    .io_a(FA_41_io_a),
    .io_b(FA_41_io_b),
    .io_cin(FA_41_io_cin)
  );
  assign io_matrix_0_0 = HA_io_s; // @[RA_Mul.scala 22:7:@1478.4]
  assign io_matrix_0_1 = io_PP_0[1]; // @[RA_Mul.scala 186:19:@1486.4]
  assign io_matrix_0_2 = FA_io_s; // @[RA_Mul.scala 47:7:@1500.4]
  assign io_matrix_0_3 = io_PP_0[3]; // @[RA_Mul.scala 192:19:@1508.4]
  assign io_matrix_0_4 = FA_1_io_s; // @[RA_Mul.scala 47:7:@1523.4]
  assign io_matrix_0_5 = FA_2_io_s; // @[RA_Mul.scala 47:7:@1540.4]
  assign io_matrix_0_6 = FA_3_io_s; // @[RA_Mul.scala 47:7:@1555.4]
  assign io_matrix_0_7 = FA_4_io_s; // @[RA_Mul.scala 47:7:@1572.4]
  assign io_matrix_0_8 = FA_5_io_s; // @[RA_Mul.scala 47:7:@1588.4]
  assign io_matrix_0_9 = FA_7_io_s; // @[RA_Mul.scala 47:7:@1613.4]
  assign io_matrix_0_10 = FA_8_io_s; // @[RA_Mul.scala 47:7:@1629.4]
  assign io_matrix_0_11 = FA_10_io_s; // @[RA_Mul.scala 47:7:@1655.4]
  assign io_matrix_0_12 = FA_12_io_s; // @[RA_Mul.scala 47:7:@1679.4]
  assign io_matrix_0_13 = FA_14_io_s; // @[RA_Mul.scala 47:7:@1705.4]
  assign io_matrix_0_14 = FA_16_io_s; // @[RA_Mul.scala 47:7:@1730.4]
  assign io_matrix_0_15 = FA_19_io_s; // @[RA_Mul.scala 47:7:@1764.4]
  assign io_matrix_0_16 = FA_21_io_s; // @[RA_Mul.scala 47:7:@1795.4]
  assign io_matrix_0_17 = FA_24_io_s; // @[RA_Mul.scala 47:7:@1828.4]
  assign io_matrix_0_18 = FA_26_io_s; // @[RA_Mul.scala 47:7:@1859.4]
  assign io_matrix_0_19 = FA_28_io_s; // @[RA_Mul.scala 47:7:@1890.4]
  assign io_matrix_0_20 = FA_30_io_s; // @[RA_Mul.scala 47:7:@1914.4]
  assign io_matrix_0_21 = FA_32_io_s; // @[RA_Mul.scala 47:7:@1939.4]
  assign io_matrix_0_22 = FA_34_io_s; // @[RA_Mul.scala 47:7:@1963.4]
  assign io_matrix_0_23 = FA_36_io_s; // @[RA_Mul.scala 47:7:@1987.4]
  assign io_matrix_0_24 = FA_37_io_s; // @[RA_Mul.scala 47:7:@2003.4]
  assign io_matrix_0_25 = FA_38_io_s; // @[RA_Mul.scala 47:7:@2020.4]
  assign io_matrix_0_26 = FA_39_io_s; // @[RA_Mul.scala 47:7:@2036.4]
  assign io_matrix_0_27 = FA_40_io_s; // @[RA_Mul.scala 47:7:@2052.4]
  assign io_matrix_0_28 = FA_41_io_s; // @[RA_Mul.scala 47:7:@2067.4]
  assign io_matrix_0_29 = io_PP_7[15]; // @[RA_Mul.scala 306:20:@2074.4]
  assign io_matrix_0_30 = io_SC[7]; // @[RA_Mul.scala 310:20:@2081.4]
  assign io_matrix_0_31 = io_SS[15]; // @[RA_Mul.scala 314:20:@2089.4]
  assign io_matrix_1_1 = HA_io_cout; // @[RA_Mul.scala 23:10:@1479.4]
  assign io_matrix_1_3 = FA_io_cout; // @[RA_Mul.scala 48:10:@1501.4]
  assign io_matrix_1_4 = io_S[2]; // @[RA_Mul.scala 197:19:@1526.4]
  assign io_matrix_1_5 = FA_1_io_cout; // @[RA_Mul.scala 48:10:@1524.4]
  assign io_matrix_1_6 = FA_2_io_cout; // @[RA_Mul.scala 48:10:@1541.4]
  assign io_matrix_1_7 = FA_3_io_cout; // @[RA_Mul.scala 48:10:@1556.4]
  assign io_matrix_1_8 = FA_4_io_cout; // @[RA_Mul.scala 48:10:@1573.4]
  assign io_matrix_1_9 = FA_5_io_cout; // @[RA_Mul.scala 48:10:@1589.4]
  assign io_matrix_1_10 = FA_7_io_cout; // @[RA_Mul.scala 48:10:@1614.4]
  assign io_matrix_1_11 = FA_8_io_cout; // @[RA_Mul.scala 48:10:@1630.4]
  assign io_matrix_1_12 = FA_10_io_cout; // @[RA_Mul.scala 48:10:@1656.4]
  assign io_matrix_1_13 = FA_12_io_cout; // @[RA_Mul.scala 48:10:@1680.4]
  assign io_matrix_1_14 = FA_14_io_cout; // @[RA_Mul.scala 48:10:@1706.4]
  assign io_matrix_1_15 = FA_16_io_cout; // @[RA_Mul.scala 48:10:@1731.4]
  assign io_matrix_1_16 = FA_19_io_cout; // @[RA_Mul.scala 48:10:@1765.4]
  assign io_matrix_1_17 = FA_21_io_cout; // @[RA_Mul.scala 48:10:@1796.4]
  assign io_matrix_1_18 = FA_24_io_cout; // @[RA_Mul.scala 48:10:@1829.4]
  assign io_matrix_1_19 = FA_26_io_cout; // @[RA_Mul.scala 48:10:@1860.4]
  assign io_matrix_1_20 = FA_28_io_cout; // @[RA_Mul.scala 48:10:@1891.4]
  assign io_matrix_1_21 = FA_30_io_cout; // @[RA_Mul.scala 48:10:@1915.4]
  assign io_matrix_1_22 = FA_32_io_cout; // @[RA_Mul.scala 48:10:@1940.4]
  assign io_matrix_1_23 = FA_34_io_cout; // @[RA_Mul.scala 48:10:@1964.4]
  assign io_matrix_1_24 = FA_36_io_cout; // @[RA_Mul.scala 48:10:@1988.4]
  assign io_matrix_1_25 = FA_37_io_cout; // @[RA_Mul.scala 48:10:@2004.4]
  assign io_matrix_1_26 = FA_38_io_cout; // @[RA_Mul.scala 48:10:@2021.4]
  assign io_matrix_1_27 = FA_39_io_cout; // @[RA_Mul.scala 48:10:@2037.4]
  assign io_matrix_1_28 = FA_40_io_cout; // @[RA_Mul.scala 48:10:@2053.4]
  assign io_matrix_1_29 = FA_41_io_cout; // @[RA_Mul.scala 48:10:@2068.4]
  assign io_matrix_1_30 = io_SS[14]; // @[RA_Mul.scala 311:20:@2083.4]
  assign io_matrix_2_3 = io_PP_1[1]; // @[RA_Mul.scala 193:19:@1510.4]
  assign io_matrix_2_6 = io_PP_3[0]; // @[RA_Mul.scala 204:19:@1558.4]
  assign io_matrix_2_7 = io_PP_3[1]; // @[RA_Mul.scala 209:19:@1575.4]
  assign io_matrix_2_8 = FA_6_io_s; // @[RA_Mul.scala 47:7:@1599.4]
  assign io_matrix_2_9 = io_PP_3[3]; // @[RA_Mul.scala 217:19:@1616.4]
  assign io_matrix_2_10 = FA_9_io_s; // @[RA_Mul.scala 47:7:@1640.4]
  assign io_matrix_2_11 = FA_11_io_s; // @[RA_Mul.scala 47:7:@1666.4]
  assign io_matrix_2_12 = FA_13_io_s; // @[RA_Mul.scala 47:7:@1690.4]
  assign io_matrix_2_13 = FA_15_io_s; // @[RA_Mul.scala 47:7:@1716.4]
  assign io_matrix_2_14 = FA_17_io_s; // @[RA_Mul.scala 47:7:@1741.4]
  assign io_matrix_2_15 = FA_20_io_s; // @[RA_Mul.scala 47:7:@1775.4]
  assign io_matrix_2_16 = FA_22_io_s; // @[RA_Mul.scala 47:7:@1806.4]
  assign io_matrix_2_17 = FA_25_io_s; // @[RA_Mul.scala 47:7:@1839.4]
  assign io_matrix_2_18 = FA_27_io_s; // @[RA_Mul.scala 47:7:@1870.4]
  assign io_matrix_2_19 = FA_29_io_s; // @[RA_Mul.scala 47:7:@1901.4]
  assign io_matrix_2_20 = FA_31_io_s; // @[RA_Mul.scala 47:7:@1925.4]
  assign io_matrix_2_21 = FA_33_io_s; // @[RA_Mul.scala 47:7:@1950.4]
  assign io_matrix_2_22 = FA_35_io_s; // @[RA_Mul.scala 47:7:@1974.4]
  assign io_matrix_2_23 = io_PP_7[9]; // @[RA_Mul.scala 283:20:@1990.4]
  assign io_matrix_2_24 = io_PP_7[10]; // @[RA_Mul.scala 288:20:@2006.4]
  assign io_matrix_2_25 = io_SS[9]; // @[RA_Mul.scala 293:20:@2023.4]
  assign io_matrix_2_26 = io_SS[10]; // @[RA_Mul.scala 297:20:@2039.4]
  assign io_matrix_2_29 = io_SS[13]; // @[RA_Mul.scala 307:20:@2076.4]
  assign io_matrix_3_6 = io_S[3]; // @[RA_Mul.scala 205:19:@1560.4]
  assign io_matrix_3_9 = FA_6_io_cout; // @[RA_Mul.scala 48:10:@1600.4]
  assign io_matrix_3_10 = io_S[5]; // @[RA_Mul.scala 223:20:@1643.4]
  assign io_matrix_3_11 = FA_9_io_cout; // @[RA_Mul.scala 48:10:@1641.4]
  assign io_matrix_3_12 = FA_11_io_cout; // @[RA_Mul.scala 48:10:@1667.4]
  assign io_matrix_3_13 = FA_13_io_cout; // @[RA_Mul.scala 48:10:@1691.4]
  assign io_matrix_3_14 = FA_15_io_cout; // @[RA_Mul.scala 48:10:@1717.4]
  assign io_matrix_3_15 = FA_17_io_cout; // @[RA_Mul.scala 48:10:@1742.4]
  assign io_matrix_3_16 = FA_20_io_cout; // @[RA_Mul.scala 48:10:@1776.4]
  assign io_matrix_3_17 = FA_22_io_cout; // @[RA_Mul.scala 48:10:@1807.4]
  assign io_matrix_3_18 = FA_25_io_cout; // @[RA_Mul.scala 48:10:@1840.4]
  assign io_matrix_3_19 = FA_27_io_cout; // @[RA_Mul.scala 48:10:@1871.4]
  assign io_matrix_3_20 = FA_29_io_cout; // @[RA_Mul.scala 48:10:@1902.4]
  assign io_matrix_3_21 = FA_31_io_cout; // @[RA_Mul.scala 48:10:@1926.4]
  assign io_matrix_3_22 = FA_33_io_cout; // @[RA_Mul.scala 48:10:@1951.4]
  assign io_matrix_3_23 = FA_35_io_cout; // @[RA_Mul.scala 48:10:@1975.4]
  assign io_matrix_3_24 = io_SS[8]; // @[RA_Mul.scala 289:20:@2008.4]
  assign io_matrix_4_9 = io_PP_4[1]; // @[RA_Mul.scala 218:19:@1618.4]
  assign io_matrix_4_12 = io_PP_6[0]; // @[RA_Mul.scala 232:20:@1693.4]
  assign io_matrix_4_13 = io_PP_6[1]; // @[RA_Mul.scala 238:20:@1719.4]
  assign io_matrix_4_14 = FA_18_io_s; // @[RA_Mul.scala 47:7:@1752.4]
  assign io_matrix_4_15 = HA_1_io_s; // @[RA_Mul.scala 22:7:@1784.4]
  assign io_matrix_4_16 = FA_23_io_s; // @[RA_Mul.scala 47:7:@1817.4]
  assign io_matrix_4_17 = HA_2_io_s; // @[RA_Mul.scala 22:7:@1848.4]
  assign io_matrix_4_18 = HA_3_io_s; // @[RA_Mul.scala 22:7:@1879.4]
  assign io_matrix_4_19 = io_SS[3]; // @[RA_Mul.scala 267:20:@1904.4]
  assign io_matrix_4_20 = io_SS[4]; // @[RA_Mul.scala 271:20:@1928.4]
  assign io_matrix_4_23 = io_SS[7]; // @[RA_Mul.scala 284:20:@1992.4]
  assign io_matrix_5_12 = io_S[6]; // @[RA_Mul.scala 233:20:@1695.4]
  assign io_matrix_5_15 = FA_18_io_cout; // @[RA_Mul.scala 48:10:@1753.4]
  assign io_matrix_5_16 = HA_1_io_cout; // @[RA_Mul.scala 23:10:@1785.4]
  assign io_matrix_5_17 = FA_23_io_cout; // @[RA_Mul.scala 48:10:@1818.4]
  assign io_matrix_5_18 = HA_2_io_cout; // @[RA_Mul.scala 23:10:@1849.4]
  assign io_matrix_5_19 = HA_3_io_cout; // @[RA_Mul.scala 23:10:@1880.4]
  assign HA_io_a = io_PP_0[0]; // @[RA_Mul.scala 20:14:@1476.4]
  assign HA_io_b = io_S[0]; // @[RA_Mul.scala 21:14:@1477.4]
  assign FA_io_a = io_PP_0[2]; // @[RA_Mul.scala 44:14:@1497.4]
  assign FA_io_b = io_PP_1[0]; // @[RA_Mul.scala 45:14:@1498.4]
  assign FA_io_cin = io_S[1]; // @[RA_Mul.scala 46:16:@1499.4]
  assign FA_1_io_a = io_PP_0[4]; // @[RA_Mul.scala 44:14:@1520.4]
  assign FA_1_io_b = io_PP_1[2]; // @[RA_Mul.scala 45:14:@1521.4]
  assign FA_1_io_cin = io_PP_2[0]; // @[RA_Mul.scala 46:16:@1522.4]
  assign FA_2_io_a = io_PP_0[5]; // @[RA_Mul.scala 44:14:@1537.4]
  assign FA_2_io_b = io_PP_1[3]; // @[RA_Mul.scala 45:14:@1538.4]
  assign FA_2_io_cin = io_PP_2[1]; // @[RA_Mul.scala 46:16:@1539.4]
  assign FA_3_io_a = io_PP_0[6]; // @[RA_Mul.scala 44:14:@1552.4]
  assign FA_3_io_b = io_PP_1[4]; // @[RA_Mul.scala 45:14:@1553.4]
  assign FA_3_io_cin = io_PP_2[2]; // @[RA_Mul.scala 46:16:@1554.4]
  assign FA_4_io_a = io_PP_0[7]; // @[RA_Mul.scala 44:14:@1569.4]
  assign FA_4_io_b = io_PP_1[5]; // @[RA_Mul.scala 45:14:@1570.4]
  assign FA_4_io_cin = io_PP_2[3]; // @[RA_Mul.scala 46:16:@1571.4]
  assign FA_5_io_a = io_PP_0[8]; // @[RA_Mul.scala 44:14:@1585.4]
  assign FA_5_io_b = io_PP_1[6]; // @[RA_Mul.scala 45:14:@1586.4]
  assign FA_5_io_cin = io_PP_2[4]; // @[RA_Mul.scala 46:16:@1587.4]
  assign FA_6_io_a = io_PP_3[2]; // @[RA_Mul.scala 44:14:@1596.4]
  assign FA_6_io_b = io_PP_4[0]; // @[RA_Mul.scala 45:14:@1597.4]
  assign FA_6_io_cin = io_S[4]; // @[RA_Mul.scala 46:16:@1598.4]
  assign FA_7_io_a = io_PP_0[9]; // @[RA_Mul.scala 44:14:@1610.4]
  assign FA_7_io_b = io_PP_1[7]; // @[RA_Mul.scala 45:14:@1611.4]
  assign FA_7_io_cin = io_PP_2[5]; // @[RA_Mul.scala 46:16:@1612.4]
  assign FA_8_io_a = io_PP_0[10]; // @[RA_Mul.scala 44:14:@1626.4]
  assign FA_8_io_b = io_PP_1[8]; // @[RA_Mul.scala 45:14:@1627.4]
  assign FA_8_io_cin = io_PP_2[6]; // @[RA_Mul.scala 46:16:@1628.4]
  assign FA_9_io_a = io_PP_3[4]; // @[RA_Mul.scala 44:14:@1637.4]
  assign FA_9_io_b = io_PP_4[2]; // @[RA_Mul.scala 45:14:@1638.4]
  assign FA_9_io_cin = io_PP_5[0]; // @[RA_Mul.scala 46:16:@1639.4]
  assign FA_10_io_a = io_PP_0[11]; // @[RA_Mul.scala 44:14:@1652.4]
  assign FA_10_io_b = io_PP_1[9]; // @[RA_Mul.scala 45:14:@1653.4]
  assign FA_10_io_cin = io_PP_2[7]; // @[RA_Mul.scala 46:16:@1654.4]
  assign FA_11_io_a = io_PP_3[5]; // @[RA_Mul.scala 44:14:@1663.4]
  assign FA_11_io_b = io_PP_4[3]; // @[RA_Mul.scala 45:14:@1664.4]
  assign FA_11_io_cin = io_PP_5[1]; // @[RA_Mul.scala 46:16:@1665.4]
  assign FA_12_io_a = io_PP_0[12]; // @[RA_Mul.scala 44:14:@1676.4]
  assign FA_12_io_b = io_PP_1[10]; // @[RA_Mul.scala 45:14:@1677.4]
  assign FA_12_io_cin = io_PP_2[8]; // @[RA_Mul.scala 46:16:@1678.4]
  assign FA_13_io_a = io_PP_3[6]; // @[RA_Mul.scala 44:14:@1687.4]
  assign FA_13_io_b = io_PP_4[4]; // @[RA_Mul.scala 45:14:@1688.4]
  assign FA_13_io_cin = io_PP_5[2]; // @[RA_Mul.scala 46:16:@1689.4]
  assign FA_14_io_a = io_PP_0[13]; // @[RA_Mul.scala 44:14:@1702.4]
  assign FA_14_io_b = io_PP_1[11]; // @[RA_Mul.scala 45:14:@1703.4]
  assign FA_14_io_cin = io_PP_2[9]; // @[RA_Mul.scala 46:16:@1704.4]
  assign FA_15_io_a = io_PP_3[7]; // @[RA_Mul.scala 44:14:@1713.4]
  assign FA_15_io_b = io_PP_4[5]; // @[RA_Mul.scala 45:14:@1714.4]
  assign FA_15_io_cin = io_PP_5[3]; // @[RA_Mul.scala 46:16:@1715.4]
  assign FA_16_io_a = io_PP_0[14]; // @[RA_Mul.scala 44:14:@1727.4]
  assign FA_16_io_b = io_PP_1[12]; // @[RA_Mul.scala 45:14:@1728.4]
  assign FA_16_io_cin = io_PP_2[10]; // @[RA_Mul.scala 46:16:@1729.4]
  assign FA_17_io_a = io_PP_3[8]; // @[RA_Mul.scala 44:14:@1738.4]
  assign FA_17_io_b = io_PP_4[6]; // @[RA_Mul.scala 45:14:@1739.4]
  assign FA_17_io_cin = io_PP_5[4]; // @[RA_Mul.scala 46:16:@1740.4]
  assign FA_18_io_a = io_PP_6[2]; // @[RA_Mul.scala 44:14:@1749.4]
  assign FA_18_io_b = io_PP_7[0]; // @[RA_Mul.scala 45:14:@1750.4]
  assign FA_18_io_cin = io_S[7]; // @[RA_Mul.scala 46:16:@1751.4]
  assign FA_19_io_a = io_PP_0[15]; // @[RA_Mul.scala 44:14:@1761.4]
  assign FA_19_io_b = io_PP_1[13]; // @[RA_Mul.scala 45:14:@1762.4]
  assign FA_19_io_cin = io_PP_2[11]; // @[RA_Mul.scala 46:16:@1763.4]
  assign FA_20_io_a = io_PP_3[9]; // @[RA_Mul.scala 44:14:@1772.4]
  assign FA_20_io_b = io_PP_4[7]; // @[RA_Mul.scala 45:14:@1773.4]
  assign FA_20_io_cin = io_PP_5[5]; // @[RA_Mul.scala 46:16:@1774.4]
  assign HA_1_io_a = io_PP_6[3]; // @[RA_Mul.scala 20:14:@1782.4]
  assign HA_1_io_b = io_PP_7[1]; // @[RA_Mul.scala 21:14:@1783.4]
  assign FA_21_io_a = io_SC[0]; // @[RA_Mul.scala 44:14:@1792.4]
  assign FA_21_io_b = io_PP_1[14]; // @[RA_Mul.scala 45:14:@1793.4]
  assign FA_21_io_cin = io_PP_2[12]; // @[RA_Mul.scala 46:16:@1794.4]
  assign FA_22_io_a = io_PP_3[10]; // @[RA_Mul.scala 44:14:@1803.4]
  assign FA_22_io_b = io_PP_4[8]; // @[RA_Mul.scala 45:14:@1804.4]
  assign FA_22_io_cin = io_PP_5[6]; // @[RA_Mul.scala 46:16:@1805.4]
  assign FA_23_io_a = io_PP_6[4]; // @[RA_Mul.scala 44:14:@1814.4]
  assign FA_23_io_b = io_PP_7[2]; // @[RA_Mul.scala 45:14:@1815.4]
  assign FA_23_io_cin = io_SS[0]; // @[RA_Mul.scala 46:16:@1816.4]
  assign FA_24_io_a = io_PP_1[15]; // @[RA_Mul.scala 44:14:@1825.4]
  assign FA_24_io_b = io_PP_2[13]; // @[RA_Mul.scala 45:14:@1826.4]
  assign FA_24_io_cin = io_PP_3[11]; // @[RA_Mul.scala 46:16:@1827.4]
  assign FA_25_io_a = io_PP_4[9]; // @[RA_Mul.scala 44:14:@1836.4]
  assign FA_25_io_b = io_PP_5[7]; // @[RA_Mul.scala 45:14:@1837.4]
  assign FA_25_io_cin = io_PP_6[5]; // @[RA_Mul.scala 46:16:@1838.4]
  assign HA_2_io_a = io_PP_7[3]; // @[RA_Mul.scala 20:14:@1846.4]
  assign HA_2_io_b = io_SS[1]; // @[RA_Mul.scala 21:14:@1847.4]
  assign FA_26_io_a = io_SC[1]; // @[RA_Mul.scala 44:14:@1856.4]
  assign FA_26_io_b = io_PP_2[14]; // @[RA_Mul.scala 45:14:@1857.4]
  assign FA_26_io_cin = io_PP_3[12]; // @[RA_Mul.scala 46:16:@1858.4]
  assign FA_27_io_a = io_PP_4[10]; // @[RA_Mul.scala 44:14:@1867.4]
  assign FA_27_io_b = io_PP_5[8]; // @[RA_Mul.scala 45:14:@1868.4]
  assign FA_27_io_cin = io_PP_6[6]; // @[RA_Mul.scala 46:16:@1869.4]
  assign HA_3_io_a = io_PP_7[4]; // @[RA_Mul.scala 20:14:@1877.4]
  assign HA_3_io_b = io_SS[2]; // @[RA_Mul.scala 21:14:@1878.4]
  assign FA_28_io_a = io_PP_2[15]; // @[RA_Mul.scala 44:14:@1887.4]
  assign FA_28_io_b = io_PP_3[13]; // @[RA_Mul.scala 45:14:@1888.4]
  assign FA_28_io_cin = io_PP_4[11]; // @[RA_Mul.scala 46:16:@1889.4]
  assign FA_29_io_a = io_PP_5[9]; // @[RA_Mul.scala 44:14:@1898.4]
  assign FA_29_io_b = io_PP_6[7]; // @[RA_Mul.scala 45:14:@1899.4]
  assign FA_29_io_cin = io_PP_7[5]; // @[RA_Mul.scala 46:16:@1900.4]
  assign FA_30_io_a = io_SC[2]; // @[RA_Mul.scala 44:14:@1911.4]
  assign FA_30_io_b = io_PP_3[14]; // @[RA_Mul.scala 45:14:@1912.4]
  assign FA_30_io_cin = io_PP_4[12]; // @[RA_Mul.scala 46:16:@1913.4]
  assign FA_31_io_a = io_PP_5[10]; // @[RA_Mul.scala 44:14:@1922.4]
  assign FA_31_io_b = io_PP_6[8]; // @[RA_Mul.scala 45:14:@1923.4]
  assign FA_31_io_cin = io_PP_7[6]; // @[RA_Mul.scala 46:16:@1924.4]
  assign FA_32_io_a = io_PP_3[15]; // @[RA_Mul.scala 44:14:@1936.4]
  assign FA_32_io_b = io_PP_4[13]; // @[RA_Mul.scala 45:14:@1937.4]
  assign FA_32_io_cin = io_PP_5[11]; // @[RA_Mul.scala 46:16:@1938.4]
  assign FA_33_io_a = io_PP_6[9]; // @[RA_Mul.scala 44:14:@1947.4]
  assign FA_33_io_b = io_PP_7[7]; // @[RA_Mul.scala 45:14:@1948.4]
  assign FA_33_io_cin = io_SS[5]; // @[RA_Mul.scala 46:16:@1949.4]
  assign FA_34_io_a = io_SC[3]; // @[RA_Mul.scala 44:14:@1960.4]
  assign FA_34_io_b = io_PP_4[14]; // @[RA_Mul.scala 45:14:@1961.4]
  assign FA_34_io_cin = io_PP_5[12]; // @[RA_Mul.scala 46:16:@1962.4]
  assign FA_35_io_a = io_PP_6[10]; // @[RA_Mul.scala 44:14:@1971.4]
  assign FA_35_io_b = io_PP_7[8]; // @[RA_Mul.scala 45:14:@1972.4]
  assign FA_35_io_cin = io_SS[6]; // @[RA_Mul.scala 46:16:@1973.4]
  assign FA_36_io_a = io_PP_4[15]; // @[RA_Mul.scala 44:14:@1984.4]
  assign FA_36_io_b = io_PP_5[13]; // @[RA_Mul.scala 45:14:@1985.4]
  assign FA_36_io_cin = io_PP_6[11]; // @[RA_Mul.scala 46:16:@1986.4]
  assign FA_37_io_a = io_SC[4]; // @[RA_Mul.scala 44:14:@2000.4]
  assign FA_37_io_b = io_PP_5[14]; // @[RA_Mul.scala 45:14:@2001.4]
  assign FA_37_io_cin = io_PP_6[12]; // @[RA_Mul.scala 46:16:@2002.4]
  assign FA_38_io_a = io_PP_5[15]; // @[RA_Mul.scala 44:14:@2017.4]
  assign FA_38_io_b = io_PP_6[13]; // @[RA_Mul.scala 45:14:@2018.4]
  assign FA_38_io_cin = io_PP_7[11]; // @[RA_Mul.scala 46:16:@2019.4]
  assign FA_39_io_a = io_SC[5]; // @[RA_Mul.scala 44:14:@2033.4]
  assign FA_39_io_b = io_PP_6[14]; // @[RA_Mul.scala 45:14:@2034.4]
  assign FA_39_io_cin = io_PP_7[12]; // @[RA_Mul.scala 46:16:@2035.4]
  assign FA_40_io_a = io_PP_6[15]; // @[RA_Mul.scala 44:14:@2049.4]
  assign FA_40_io_b = io_PP_7[13]; // @[RA_Mul.scala 45:14:@2050.4]
  assign FA_40_io_cin = io_SS[11]; // @[RA_Mul.scala 46:16:@2051.4]
  assign FA_41_io_a = io_SC[6]; // @[RA_Mul.scala 44:14:@2064.4]
  assign FA_41_io_b = io_PP_7[14]; // @[RA_Mul.scala 45:14:@2065.4]
  assign FA_41_io_cin = io_SS[12]; // @[RA_Mul.scala 46:16:@2066.4]
endmodule
module Reduction_2( // @[:@2571.2]
  output  io_matrix_o_0_0, // @[:@2574.4]
  output  io_matrix_o_0_1, // @[:@2574.4]
  output  io_matrix_o_0_2, // @[:@2574.4]
  output  io_matrix_o_0_3, // @[:@2574.4]
  output  io_matrix_o_0_4, // @[:@2574.4]
  output  io_matrix_o_0_5, // @[:@2574.4]
  output  io_matrix_o_0_6, // @[:@2574.4]
  output  io_matrix_o_0_7, // @[:@2574.4]
  output  io_matrix_o_0_8, // @[:@2574.4]
  output  io_matrix_o_0_9, // @[:@2574.4]
  output  io_matrix_o_0_10, // @[:@2574.4]
  output  io_matrix_o_0_11, // @[:@2574.4]
  output  io_matrix_o_0_12, // @[:@2574.4]
  output  io_matrix_o_0_13, // @[:@2574.4]
  output  io_matrix_o_0_14, // @[:@2574.4]
  output  io_matrix_o_0_15, // @[:@2574.4]
  output  io_matrix_o_0_16, // @[:@2574.4]
  output  io_matrix_o_0_17, // @[:@2574.4]
  output  io_matrix_o_0_18, // @[:@2574.4]
  output  io_matrix_o_0_19, // @[:@2574.4]
  output  io_matrix_o_0_20, // @[:@2574.4]
  output  io_matrix_o_0_21, // @[:@2574.4]
  output  io_matrix_o_0_22, // @[:@2574.4]
  output  io_matrix_o_0_23, // @[:@2574.4]
  output  io_matrix_o_0_24, // @[:@2574.4]
  output  io_matrix_o_0_25, // @[:@2574.4]
  output  io_matrix_o_0_26, // @[:@2574.4]
  output  io_matrix_o_0_27, // @[:@2574.4]
  output  io_matrix_o_0_28, // @[:@2574.4]
  output  io_matrix_o_0_29, // @[:@2574.4]
  output  io_matrix_o_0_30, // @[:@2574.4]
  output  io_matrix_o_0_31, // @[:@2574.4]
  output  io_matrix_o_1_2, // @[:@2574.4]
  output  io_matrix_o_1_4, // @[:@2574.4]
  output  io_matrix_o_1_5, // @[:@2574.4]
  output  io_matrix_o_1_6, // @[:@2574.4]
  output  io_matrix_o_1_7, // @[:@2574.4]
  output  io_matrix_o_1_8, // @[:@2574.4]
  output  io_matrix_o_1_9, // @[:@2574.4]
  output  io_matrix_o_1_10, // @[:@2574.4]
  output  io_matrix_o_1_11, // @[:@2574.4]
  output  io_matrix_o_1_12, // @[:@2574.4]
  output  io_matrix_o_1_13, // @[:@2574.4]
  output  io_matrix_o_1_14, // @[:@2574.4]
  output  io_matrix_o_1_15, // @[:@2574.4]
  output  io_matrix_o_1_16, // @[:@2574.4]
  output  io_matrix_o_1_17, // @[:@2574.4]
  output  io_matrix_o_1_18, // @[:@2574.4]
  output  io_matrix_o_1_19, // @[:@2574.4]
  output  io_matrix_o_1_20, // @[:@2574.4]
  output  io_matrix_o_1_21, // @[:@2574.4]
  output  io_matrix_o_1_22, // @[:@2574.4]
  output  io_matrix_o_1_23, // @[:@2574.4]
  output  io_matrix_o_1_24, // @[:@2574.4]
  output  io_matrix_o_1_25, // @[:@2574.4]
  output  io_matrix_o_1_26, // @[:@2574.4]
  output  io_matrix_o_1_27, // @[:@2574.4]
  output  io_matrix_o_1_28, // @[:@2574.4]
  output  io_matrix_o_1_30, // @[:@2574.4]
  output  io_matrix_o_2_4, // @[:@2574.4]
  output  io_matrix_o_2_9, // @[:@2574.4]
  output  io_matrix_o_2_10, // @[:@2574.4]
  output  io_matrix_o_2_11, // @[:@2574.4]
  output  io_matrix_o_2_12, // @[:@2574.4]
  output  io_matrix_o_2_13, // @[:@2574.4]
  output  io_matrix_o_2_14, // @[:@2574.4]
  output  io_matrix_o_2_15, // @[:@2574.4]
  output  io_matrix_o_2_16, // @[:@2574.4]
  output  io_matrix_o_2_17, // @[:@2574.4]
  output  io_matrix_o_2_18, // @[:@2574.4]
  output  io_matrix_o_2_19, // @[:@2574.4]
  output  io_matrix_o_2_20, // @[:@2574.4]
  output  io_matrix_o_2_21, // @[:@2574.4]
  output  io_matrix_o_2_22, // @[:@2574.4]
  output  io_matrix_o_2_23, // @[:@2574.4]
  output  io_matrix_o_2_24, // @[:@2574.4]
  output  io_matrix_o_2_27, // @[:@2574.4]
  output  io_matrix_o_2_30, // @[:@2574.4]
  output  io_matrix_o_3_9, // @[:@2574.4]
  output  io_matrix_o_3_13, // @[:@2574.4]
  output  io_matrix_o_3_14, // @[:@2574.4]
  output  io_matrix_o_3_15, // @[:@2574.4]
  output  io_matrix_o_3_16, // @[:@2574.4]
  output  io_matrix_o_3_17, // @[:@2574.4]
  output  io_matrix_o_3_18, // @[:@2574.4]
  output  io_matrix_o_3_19, // @[:@2574.4]
  output  io_matrix_o_3_20, // @[:@2574.4]
  output  io_matrix_o_3_21, // @[:@2574.4]
  output  io_matrix_o_3_23, // @[:@2574.4]
  input   io_matrix_i_0_0, // @[:@2574.4]
  input   io_matrix_i_0_1, // @[:@2574.4]
  input   io_matrix_i_0_2, // @[:@2574.4]
  input   io_matrix_i_0_3, // @[:@2574.4]
  input   io_matrix_i_0_4, // @[:@2574.4]
  input   io_matrix_i_0_5, // @[:@2574.4]
  input   io_matrix_i_0_6, // @[:@2574.4]
  input   io_matrix_i_0_7, // @[:@2574.4]
  input   io_matrix_i_0_8, // @[:@2574.4]
  input   io_matrix_i_0_9, // @[:@2574.4]
  input   io_matrix_i_0_10, // @[:@2574.4]
  input   io_matrix_i_0_11, // @[:@2574.4]
  input   io_matrix_i_0_12, // @[:@2574.4]
  input   io_matrix_i_0_13, // @[:@2574.4]
  input   io_matrix_i_0_14, // @[:@2574.4]
  input   io_matrix_i_0_15, // @[:@2574.4]
  input   io_matrix_i_0_16, // @[:@2574.4]
  input   io_matrix_i_0_17, // @[:@2574.4]
  input   io_matrix_i_0_18, // @[:@2574.4]
  input   io_matrix_i_0_19, // @[:@2574.4]
  input   io_matrix_i_0_20, // @[:@2574.4]
  input   io_matrix_i_0_21, // @[:@2574.4]
  input   io_matrix_i_0_22, // @[:@2574.4]
  input   io_matrix_i_0_23, // @[:@2574.4]
  input   io_matrix_i_0_24, // @[:@2574.4]
  input   io_matrix_i_0_25, // @[:@2574.4]
  input   io_matrix_i_0_26, // @[:@2574.4]
  input   io_matrix_i_0_27, // @[:@2574.4]
  input   io_matrix_i_0_28, // @[:@2574.4]
  input   io_matrix_i_0_29, // @[:@2574.4]
  input   io_matrix_i_0_30, // @[:@2574.4]
  input   io_matrix_i_0_31, // @[:@2574.4]
  input   io_matrix_i_1_1, // @[:@2574.4]
  input   io_matrix_i_1_3, // @[:@2574.4]
  input   io_matrix_i_1_4, // @[:@2574.4]
  input   io_matrix_i_1_5, // @[:@2574.4]
  input   io_matrix_i_1_6, // @[:@2574.4]
  input   io_matrix_i_1_7, // @[:@2574.4]
  input   io_matrix_i_1_8, // @[:@2574.4]
  input   io_matrix_i_1_9, // @[:@2574.4]
  input   io_matrix_i_1_10, // @[:@2574.4]
  input   io_matrix_i_1_11, // @[:@2574.4]
  input   io_matrix_i_1_12, // @[:@2574.4]
  input   io_matrix_i_1_13, // @[:@2574.4]
  input   io_matrix_i_1_14, // @[:@2574.4]
  input   io_matrix_i_1_15, // @[:@2574.4]
  input   io_matrix_i_1_16, // @[:@2574.4]
  input   io_matrix_i_1_17, // @[:@2574.4]
  input   io_matrix_i_1_18, // @[:@2574.4]
  input   io_matrix_i_1_19, // @[:@2574.4]
  input   io_matrix_i_1_20, // @[:@2574.4]
  input   io_matrix_i_1_21, // @[:@2574.4]
  input   io_matrix_i_1_22, // @[:@2574.4]
  input   io_matrix_i_1_23, // @[:@2574.4]
  input   io_matrix_i_1_24, // @[:@2574.4]
  input   io_matrix_i_1_25, // @[:@2574.4]
  input   io_matrix_i_1_26, // @[:@2574.4]
  input   io_matrix_i_1_27, // @[:@2574.4]
  input   io_matrix_i_1_28, // @[:@2574.4]
  input   io_matrix_i_1_29, // @[:@2574.4]
  input   io_matrix_i_1_30, // @[:@2574.4]
  input   io_matrix_i_2_3, // @[:@2574.4]
  input   io_matrix_i_2_6, // @[:@2574.4]
  input   io_matrix_i_2_7, // @[:@2574.4]
  input   io_matrix_i_2_8, // @[:@2574.4]
  input   io_matrix_i_2_9, // @[:@2574.4]
  input   io_matrix_i_2_10, // @[:@2574.4]
  input   io_matrix_i_2_11, // @[:@2574.4]
  input   io_matrix_i_2_12, // @[:@2574.4]
  input   io_matrix_i_2_13, // @[:@2574.4]
  input   io_matrix_i_2_14, // @[:@2574.4]
  input   io_matrix_i_2_15, // @[:@2574.4]
  input   io_matrix_i_2_16, // @[:@2574.4]
  input   io_matrix_i_2_17, // @[:@2574.4]
  input   io_matrix_i_2_18, // @[:@2574.4]
  input   io_matrix_i_2_19, // @[:@2574.4]
  input   io_matrix_i_2_20, // @[:@2574.4]
  input   io_matrix_i_2_21, // @[:@2574.4]
  input   io_matrix_i_2_22, // @[:@2574.4]
  input   io_matrix_i_2_23, // @[:@2574.4]
  input   io_matrix_i_2_24, // @[:@2574.4]
  input   io_matrix_i_2_25, // @[:@2574.4]
  input   io_matrix_i_2_26, // @[:@2574.4]
  input   io_matrix_i_2_29, // @[:@2574.4]
  input   io_matrix_i_3_6, // @[:@2574.4]
  input   io_matrix_i_3_9, // @[:@2574.4]
  input   io_matrix_i_3_10, // @[:@2574.4]
  input   io_matrix_i_3_11, // @[:@2574.4]
  input   io_matrix_i_3_12, // @[:@2574.4]
  input   io_matrix_i_3_13, // @[:@2574.4]
  input   io_matrix_i_3_14, // @[:@2574.4]
  input   io_matrix_i_3_15, // @[:@2574.4]
  input   io_matrix_i_3_16, // @[:@2574.4]
  input   io_matrix_i_3_17, // @[:@2574.4]
  input   io_matrix_i_3_18, // @[:@2574.4]
  input   io_matrix_i_3_19, // @[:@2574.4]
  input   io_matrix_i_3_20, // @[:@2574.4]
  input   io_matrix_i_3_21, // @[:@2574.4]
  input   io_matrix_i_3_22, // @[:@2574.4]
  input   io_matrix_i_3_23, // @[:@2574.4]
  input   io_matrix_i_3_24, // @[:@2574.4]
  input   io_matrix_i_4_9, // @[:@2574.4]
  input   io_matrix_i_4_12, // @[:@2574.4]
  input   io_matrix_i_4_13, // @[:@2574.4]
  input   io_matrix_i_4_14, // @[:@2574.4]
  input   io_matrix_i_4_15, // @[:@2574.4]
  input   io_matrix_i_4_16, // @[:@2574.4]
  input   io_matrix_i_4_17, // @[:@2574.4]
  input   io_matrix_i_4_18, // @[:@2574.4]
  input   io_matrix_i_4_19, // @[:@2574.4]
  input   io_matrix_i_4_20, // @[:@2574.4]
  input   io_matrix_i_4_23, // @[:@2574.4]
  input   io_matrix_i_5_12, // @[:@2574.4]
  input   io_matrix_i_5_15, // @[:@2574.4]
  input   io_matrix_i_5_16, // @[:@2574.4]
  input   io_matrix_i_5_17, // @[:@2574.4]
  input   io_matrix_i_5_18, // @[:@2574.4]
  input   io_matrix_i_5_19 // @[:@2574.4]
);
  wire  HA_io_s; // @[RA_Mul.scala 19:21:@2580.4]
  wire  HA_io_cout; // @[RA_Mul.scala 19:21:@2580.4]
  wire  HA_io_a; // @[RA_Mul.scala 19:21:@2580.4]
  wire  HA_io_b; // @[RA_Mul.scala 19:21:@2580.4]
  wire  FA_io_s; // @[RA_Mul.scala 43:21:@2593.4]
  wire  FA_io_cout; // @[RA_Mul.scala 43:21:@2593.4]
  wire  FA_io_a; // @[RA_Mul.scala 43:21:@2593.4]
  wire  FA_io_b; // @[RA_Mul.scala 43:21:@2593.4]
  wire  FA_io_cin; // @[RA_Mul.scala 43:21:@2593.4]
  wire  FA_1_io_s; // @[RA_Mul.scala 43:21:@2611.4]
  wire  FA_1_io_cout; // @[RA_Mul.scala 43:21:@2611.4]
  wire  FA_1_io_a; // @[RA_Mul.scala 43:21:@2611.4]
  wire  FA_1_io_b; // @[RA_Mul.scala 43:21:@2611.4]
  wire  FA_1_io_cin; // @[RA_Mul.scala 43:21:@2611.4]
  wire  FA_2_io_s; // @[RA_Mul.scala 43:21:@2622.4]
  wire  FA_2_io_cout; // @[RA_Mul.scala 43:21:@2622.4]
  wire  FA_2_io_a; // @[RA_Mul.scala 43:21:@2622.4]
  wire  FA_2_io_b; // @[RA_Mul.scala 43:21:@2622.4]
  wire  FA_2_io_cin; // @[RA_Mul.scala 43:21:@2622.4]
  wire  FA_3_io_s; // @[RA_Mul.scala 43:21:@2632.4]
  wire  FA_3_io_cout; // @[RA_Mul.scala 43:21:@2632.4]
  wire  FA_3_io_a; // @[RA_Mul.scala 43:21:@2632.4]
  wire  FA_3_io_b; // @[RA_Mul.scala 43:21:@2632.4]
  wire  FA_3_io_cin; // @[RA_Mul.scala 43:21:@2632.4]
  wire  FA_4_io_s; // @[RA_Mul.scala 43:21:@2642.4]
  wire  FA_4_io_cout; // @[RA_Mul.scala 43:21:@2642.4]
  wire  FA_4_io_a; // @[RA_Mul.scala 43:21:@2642.4]
  wire  FA_4_io_b; // @[RA_Mul.scala 43:21:@2642.4]
  wire  FA_4_io_cin; // @[RA_Mul.scala 43:21:@2642.4]
  wire  FA_5_io_s; // @[RA_Mul.scala 43:21:@2652.4]
  wire  FA_5_io_cout; // @[RA_Mul.scala 43:21:@2652.4]
  wire  FA_5_io_a; // @[RA_Mul.scala 43:21:@2652.4]
  wire  FA_5_io_b; // @[RA_Mul.scala 43:21:@2652.4]
  wire  FA_5_io_cin; // @[RA_Mul.scala 43:21:@2652.4]
  wire  FA_6_io_s; // @[RA_Mul.scala 43:21:@2662.4]
  wire  FA_6_io_cout; // @[RA_Mul.scala 43:21:@2662.4]
  wire  FA_6_io_a; // @[RA_Mul.scala 43:21:@2662.4]
  wire  FA_6_io_b; // @[RA_Mul.scala 43:21:@2662.4]
  wire  FA_6_io_cin; // @[RA_Mul.scala 43:21:@2662.4]
  wire  FA_7_io_s; // @[RA_Mul.scala 43:21:@2672.4]
  wire  FA_7_io_cout; // @[RA_Mul.scala 43:21:@2672.4]
  wire  FA_7_io_a; // @[RA_Mul.scala 43:21:@2672.4]
  wire  FA_7_io_b; // @[RA_Mul.scala 43:21:@2672.4]
  wire  FA_7_io_cin; // @[RA_Mul.scala 43:21:@2672.4]
  wire  FA_8_io_s; // @[RA_Mul.scala 43:21:@2680.4]
  wire  FA_8_io_cout; // @[RA_Mul.scala 43:21:@2680.4]
  wire  FA_8_io_a; // @[RA_Mul.scala 43:21:@2680.4]
  wire  FA_8_io_b; // @[RA_Mul.scala 43:21:@2680.4]
  wire  FA_8_io_cin; // @[RA_Mul.scala 43:21:@2680.4]
  wire  FA_9_io_s; // @[RA_Mul.scala 43:21:@2689.4]
  wire  FA_9_io_cout; // @[RA_Mul.scala 43:21:@2689.4]
  wire  FA_9_io_a; // @[RA_Mul.scala 43:21:@2689.4]
  wire  FA_9_io_b; // @[RA_Mul.scala 43:21:@2689.4]
  wire  FA_9_io_cin; // @[RA_Mul.scala 43:21:@2689.4]
  wire  HA_1_io_s; // @[RA_Mul.scala 19:21:@2697.4]
  wire  HA_1_io_cout; // @[RA_Mul.scala 19:21:@2697.4]
  wire  HA_1_io_a; // @[RA_Mul.scala 19:21:@2697.4]
  wire  HA_1_io_b; // @[RA_Mul.scala 19:21:@2697.4]
  wire  FA_10_io_s; // @[RA_Mul.scala 43:21:@2704.4]
  wire  FA_10_io_cout; // @[RA_Mul.scala 43:21:@2704.4]
  wire  FA_10_io_a; // @[RA_Mul.scala 43:21:@2704.4]
  wire  FA_10_io_b; // @[RA_Mul.scala 43:21:@2704.4]
  wire  FA_10_io_cin; // @[RA_Mul.scala 43:21:@2704.4]
  wire  HA_2_io_s; // @[RA_Mul.scala 19:21:@2712.4]
  wire  HA_2_io_cout; // @[RA_Mul.scala 19:21:@2712.4]
  wire  HA_2_io_a; // @[RA_Mul.scala 19:21:@2712.4]
  wire  HA_2_io_b; // @[RA_Mul.scala 19:21:@2712.4]
  wire  FA_11_io_s; // @[RA_Mul.scala 43:21:@2719.4]
  wire  FA_11_io_cout; // @[RA_Mul.scala 43:21:@2719.4]
  wire  FA_11_io_a; // @[RA_Mul.scala 43:21:@2719.4]
  wire  FA_11_io_b; // @[RA_Mul.scala 43:21:@2719.4]
  wire  FA_11_io_cin; // @[RA_Mul.scala 43:21:@2719.4]
  wire  FA_12_io_s; // @[RA_Mul.scala 43:21:@2727.4]
  wire  FA_12_io_cout; // @[RA_Mul.scala 43:21:@2727.4]
  wire  FA_12_io_a; // @[RA_Mul.scala 43:21:@2727.4]
  wire  FA_12_io_b; // @[RA_Mul.scala 43:21:@2727.4]
  wire  FA_12_io_cin; // @[RA_Mul.scala 43:21:@2727.4]
  wire  FA_13_io_s; // @[RA_Mul.scala 43:21:@2735.4]
  wire  FA_13_io_cout; // @[RA_Mul.scala 43:21:@2735.4]
  wire  FA_13_io_a; // @[RA_Mul.scala 43:21:@2735.4]
  wire  FA_13_io_b; // @[RA_Mul.scala 43:21:@2735.4]
  wire  FA_13_io_cin; // @[RA_Mul.scala 43:21:@2735.4]
  wire  FA_14_io_s; // @[RA_Mul.scala 43:21:@2743.4]
  wire  FA_14_io_cout; // @[RA_Mul.scala 43:21:@2743.4]
  wire  FA_14_io_a; // @[RA_Mul.scala 43:21:@2743.4]
  wire  FA_14_io_b; // @[RA_Mul.scala 43:21:@2743.4]
  wire  FA_14_io_cin; // @[RA_Mul.scala 43:21:@2743.4]
  wire  FA_15_io_s; // @[RA_Mul.scala 43:21:@2751.4]
  wire  FA_15_io_cout; // @[RA_Mul.scala 43:21:@2751.4]
  wire  FA_15_io_a; // @[RA_Mul.scala 43:21:@2751.4]
  wire  FA_15_io_b; // @[RA_Mul.scala 43:21:@2751.4]
  wire  FA_15_io_cin; // @[RA_Mul.scala 43:21:@2751.4]
  wire  FA_16_io_s; // @[RA_Mul.scala 43:21:@2759.4]
  wire  FA_16_io_cout; // @[RA_Mul.scala 43:21:@2759.4]
  wire  FA_16_io_a; // @[RA_Mul.scala 43:21:@2759.4]
  wire  FA_16_io_b; // @[RA_Mul.scala 43:21:@2759.4]
  wire  FA_16_io_cin; // @[RA_Mul.scala 43:21:@2759.4]
  wire  FA_17_io_s; // @[RA_Mul.scala 43:21:@2767.4]
  wire  FA_17_io_cout; // @[RA_Mul.scala 43:21:@2767.4]
  wire  FA_17_io_a; // @[RA_Mul.scala 43:21:@2767.4]
  wire  FA_17_io_b; // @[RA_Mul.scala 43:21:@2767.4]
  wire  FA_17_io_cin; // @[RA_Mul.scala 43:21:@2767.4]
  wire  FA_18_io_s; // @[RA_Mul.scala 43:21:@2775.4]
  wire  FA_18_io_cout; // @[RA_Mul.scala 43:21:@2775.4]
  wire  FA_18_io_a; // @[RA_Mul.scala 43:21:@2775.4]
  wire  FA_18_io_b; // @[RA_Mul.scala 43:21:@2775.4]
  wire  FA_18_io_cin; // @[RA_Mul.scala 43:21:@2775.4]
  wire  FA_19_io_s; // @[RA_Mul.scala 43:21:@2783.4]
  wire  FA_19_io_cout; // @[RA_Mul.scala 43:21:@2783.4]
  wire  FA_19_io_a; // @[RA_Mul.scala 43:21:@2783.4]
  wire  FA_19_io_b; // @[RA_Mul.scala 43:21:@2783.4]
  wire  FA_19_io_cin; // @[RA_Mul.scala 43:21:@2783.4]
  wire  FA_20_io_s; // @[RA_Mul.scala 43:21:@2791.4]
  wire  FA_20_io_cout; // @[RA_Mul.scala 43:21:@2791.4]
  wire  FA_20_io_a; // @[RA_Mul.scala 43:21:@2791.4]
  wire  FA_20_io_b; // @[RA_Mul.scala 43:21:@2791.4]
  wire  FA_20_io_cin; // @[RA_Mul.scala 43:21:@2791.4]
  wire  FA_21_io_s; // @[RA_Mul.scala 43:21:@2799.4]
  wire  FA_21_io_cout; // @[RA_Mul.scala 43:21:@2799.4]
  wire  FA_21_io_a; // @[RA_Mul.scala 43:21:@2799.4]
  wire  FA_21_io_b; // @[RA_Mul.scala 43:21:@2799.4]
  wire  FA_21_io_cin; // @[RA_Mul.scala 43:21:@2799.4]
  wire  HA_3_io_s; // @[RA_Mul.scala 19:21:@2807.4]
  wire  HA_3_io_cout; // @[RA_Mul.scala 19:21:@2807.4]
  wire  HA_3_io_a; // @[RA_Mul.scala 19:21:@2807.4]
  wire  HA_3_io_b; // @[RA_Mul.scala 19:21:@2807.4]
  wire  FA_22_io_s; // @[RA_Mul.scala 43:21:@2814.4]
  wire  FA_22_io_cout; // @[RA_Mul.scala 43:21:@2814.4]
  wire  FA_22_io_a; // @[RA_Mul.scala 43:21:@2814.4]
  wire  FA_22_io_b; // @[RA_Mul.scala 43:21:@2814.4]
  wire  FA_22_io_cin; // @[RA_Mul.scala 43:21:@2814.4]
  wire  FA_23_io_s; // @[RA_Mul.scala 43:21:@2823.4]
  wire  FA_23_io_cout; // @[RA_Mul.scala 43:21:@2823.4]
  wire  FA_23_io_a; // @[RA_Mul.scala 43:21:@2823.4]
  wire  FA_23_io_b; // @[RA_Mul.scala 43:21:@2823.4]
  wire  FA_23_io_cin; // @[RA_Mul.scala 43:21:@2823.4]
  wire  FA_24_io_s; // @[RA_Mul.scala 43:21:@2833.4]
  wire  FA_24_io_cout; // @[RA_Mul.scala 43:21:@2833.4]
  wire  FA_24_io_a; // @[RA_Mul.scala 43:21:@2833.4]
  wire  FA_24_io_b; // @[RA_Mul.scala 43:21:@2833.4]
  wire  FA_24_io_cin; // @[RA_Mul.scala 43:21:@2833.4]
  wire  FA_25_io_s; // @[RA_Mul.scala 43:21:@2843.4]
  wire  FA_25_io_cout; // @[RA_Mul.scala 43:21:@2843.4]
  wire  FA_25_io_a; // @[RA_Mul.scala 43:21:@2843.4]
  wire  FA_25_io_b; // @[RA_Mul.scala 43:21:@2843.4]
  wire  FA_25_io_cin; // @[RA_Mul.scala 43:21:@2843.4]
  wire  FA_26_io_s; // @[RA_Mul.scala 43:21:@2853.4]
  wire  FA_26_io_cout; // @[RA_Mul.scala 43:21:@2853.4]
  wire  FA_26_io_a; // @[RA_Mul.scala 43:21:@2853.4]
  wire  FA_26_io_b; // @[RA_Mul.scala 43:21:@2853.4]
  wire  FA_26_io_cin; // @[RA_Mul.scala 43:21:@2853.4]
  wire  FA_27_io_s; // @[RA_Mul.scala 43:21:@2863.4]
  wire  FA_27_io_cout; // @[RA_Mul.scala 43:21:@2863.4]
  wire  FA_27_io_a; // @[RA_Mul.scala 43:21:@2863.4]
  wire  FA_27_io_b; // @[RA_Mul.scala 43:21:@2863.4]
  wire  FA_27_io_cin; // @[RA_Mul.scala 43:21:@2863.4]
  wire  FA_28_io_s; // @[RA_Mul.scala 43:21:@2880.4]
  wire  FA_28_io_cout; // @[RA_Mul.scala 43:21:@2880.4]
  wire  FA_28_io_a; // @[RA_Mul.scala 43:21:@2880.4]
  wire  FA_28_io_b; // @[RA_Mul.scala 43:21:@2880.4]
  wire  FA_28_io_cin; // @[RA_Mul.scala 43:21:@2880.4]
  HA HA ( // @[RA_Mul.scala 19:21:@2580.4]
    .io_s(HA_io_s),
    .io_cout(HA_io_cout),
    .io_a(HA_io_a),
    .io_b(HA_io_b)
  );
  FA FA ( // @[RA_Mul.scala 43:21:@2593.4]
    .io_s(FA_io_s),
    .io_cout(FA_io_cout),
    .io_a(FA_io_a),
    .io_b(FA_io_b),
    .io_cin(FA_io_cin)
  );
  FA FA_1 ( // @[RA_Mul.scala 43:21:@2611.4]
    .io_s(FA_1_io_s),
    .io_cout(FA_1_io_cout),
    .io_a(FA_1_io_a),
    .io_b(FA_1_io_b),
    .io_cin(FA_1_io_cin)
  );
  FA FA_2 ( // @[RA_Mul.scala 43:21:@2622.4]
    .io_s(FA_2_io_s),
    .io_cout(FA_2_io_cout),
    .io_a(FA_2_io_a),
    .io_b(FA_2_io_b),
    .io_cin(FA_2_io_cin)
  );
  FA FA_3 ( // @[RA_Mul.scala 43:21:@2632.4]
    .io_s(FA_3_io_s),
    .io_cout(FA_3_io_cout),
    .io_a(FA_3_io_a),
    .io_b(FA_3_io_b),
    .io_cin(FA_3_io_cin)
  );
  FA FA_4 ( // @[RA_Mul.scala 43:21:@2642.4]
    .io_s(FA_4_io_s),
    .io_cout(FA_4_io_cout),
    .io_a(FA_4_io_a),
    .io_b(FA_4_io_b),
    .io_cin(FA_4_io_cin)
  );
  FA FA_5 ( // @[RA_Mul.scala 43:21:@2652.4]
    .io_s(FA_5_io_s),
    .io_cout(FA_5_io_cout),
    .io_a(FA_5_io_a),
    .io_b(FA_5_io_b),
    .io_cin(FA_5_io_cin)
  );
  FA FA_6 ( // @[RA_Mul.scala 43:21:@2662.4]
    .io_s(FA_6_io_s),
    .io_cout(FA_6_io_cout),
    .io_a(FA_6_io_a),
    .io_b(FA_6_io_b),
    .io_cin(FA_6_io_cin)
  );
  FA FA_7 ( // @[RA_Mul.scala 43:21:@2672.4]
    .io_s(FA_7_io_s),
    .io_cout(FA_7_io_cout),
    .io_a(FA_7_io_a),
    .io_b(FA_7_io_b),
    .io_cin(FA_7_io_cin)
  );
  FA FA_8 ( // @[RA_Mul.scala 43:21:@2680.4]
    .io_s(FA_8_io_s),
    .io_cout(FA_8_io_cout),
    .io_a(FA_8_io_a),
    .io_b(FA_8_io_b),
    .io_cin(FA_8_io_cin)
  );
  FA FA_9 ( // @[RA_Mul.scala 43:21:@2689.4]
    .io_s(FA_9_io_s),
    .io_cout(FA_9_io_cout),
    .io_a(FA_9_io_a),
    .io_b(FA_9_io_b),
    .io_cin(FA_9_io_cin)
  );
  HA HA_1 ( // @[RA_Mul.scala 19:21:@2697.4]
    .io_s(HA_1_io_s),
    .io_cout(HA_1_io_cout),
    .io_a(HA_1_io_a),
    .io_b(HA_1_io_b)
  );
  FA FA_10 ( // @[RA_Mul.scala 43:21:@2704.4]
    .io_s(FA_10_io_s),
    .io_cout(FA_10_io_cout),
    .io_a(FA_10_io_a),
    .io_b(FA_10_io_b),
    .io_cin(FA_10_io_cin)
  );
  HA HA_2 ( // @[RA_Mul.scala 19:21:@2712.4]
    .io_s(HA_2_io_s),
    .io_cout(HA_2_io_cout),
    .io_a(HA_2_io_a),
    .io_b(HA_2_io_b)
  );
  FA FA_11 ( // @[RA_Mul.scala 43:21:@2719.4]
    .io_s(FA_11_io_s),
    .io_cout(FA_11_io_cout),
    .io_a(FA_11_io_a),
    .io_b(FA_11_io_b),
    .io_cin(FA_11_io_cin)
  );
  FA FA_12 ( // @[RA_Mul.scala 43:21:@2727.4]
    .io_s(FA_12_io_s),
    .io_cout(FA_12_io_cout),
    .io_a(FA_12_io_a),
    .io_b(FA_12_io_b),
    .io_cin(FA_12_io_cin)
  );
  FA FA_13 ( // @[RA_Mul.scala 43:21:@2735.4]
    .io_s(FA_13_io_s),
    .io_cout(FA_13_io_cout),
    .io_a(FA_13_io_a),
    .io_b(FA_13_io_b),
    .io_cin(FA_13_io_cin)
  );
  FA FA_14 ( // @[RA_Mul.scala 43:21:@2743.4]
    .io_s(FA_14_io_s),
    .io_cout(FA_14_io_cout),
    .io_a(FA_14_io_a),
    .io_b(FA_14_io_b),
    .io_cin(FA_14_io_cin)
  );
  FA FA_15 ( // @[RA_Mul.scala 43:21:@2751.4]
    .io_s(FA_15_io_s),
    .io_cout(FA_15_io_cout),
    .io_a(FA_15_io_a),
    .io_b(FA_15_io_b),
    .io_cin(FA_15_io_cin)
  );
  FA FA_16 ( // @[RA_Mul.scala 43:21:@2759.4]
    .io_s(FA_16_io_s),
    .io_cout(FA_16_io_cout),
    .io_a(FA_16_io_a),
    .io_b(FA_16_io_b),
    .io_cin(FA_16_io_cin)
  );
  FA FA_17 ( // @[RA_Mul.scala 43:21:@2767.4]
    .io_s(FA_17_io_s),
    .io_cout(FA_17_io_cout),
    .io_a(FA_17_io_a),
    .io_b(FA_17_io_b),
    .io_cin(FA_17_io_cin)
  );
  FA FA_18 ( // @[RA_Mul.scala 43:21:@2775.4]
    .io_s(FA_18_io_s),
    .io_cout(FA_18_io_cout),
    .io_a(FA_18_io_a),
    .io_b(FA_18_io_b),
    .io_cin(FA_18_io_cin)
  );
  FA FA_19 ( // @[RA_Mul.scala 43:21:@2783.4]
    .io_s(FA_19_io_s),
    .io_cout(FA_19_io_cout),
    .io_a(FA_19_io_a),
    .io_b(FA_19_io_b),
    .io_cin(FA_19_io_cin)
  );
  FA FA_20 ( // @[RA_Mul.scala 43:21:@2791.4]
    .io_s(FA_20_io_s),
    .io_cout(FA_20_io_cout),
    .io_a(FA_20_io_a),
    .io_b(FA_20_io_b),
    .io_cin(FA_20_io_cin)
  );
  FA FA_21 ( // @[RA_Mul.scala 43:21:@2799.4]
    .io_s(FA_21_io_s),
    .io_cout(FA_21_io_cout),
    .io_a(FA_21_io_a),
    .io_b(FA_21_io_b),
    .io_cin(FA_21_io_cin)
  );
  HA HA_3 ( // @[RA_Mul.scala 19:21:@2807.4]
    .io_s(HA_3_io_s),
    .io_cout(HA_3_io_cout),
    .io_a(HA_3_io_a),
    .io_b(HA_3_io_b)
  );
  FA FA_22 ( // @[RA_Mul.scala 43:21:@2814.4]
    .io_s(FA_22_io_s),
    .io_cout(FA_22_io_cout),
    .io_a(FA_22_io_a),
    .io_b(FA_22_io_b),
    .io_cin(FA_22_io_cin)
  );
  FA FA_23 ( // @[RA_Mul.scala 43:21:@2823.4]
    .io_s(FA_23_io_s),
    .io_cout(FA_23_io_cout),
    .io_a(FA_23_io_a),
    .io_b(FA_23_io_b),
    .io_cin(FA_23_io_cin)
  );
  FA FA_24 ( // @[RA_Mul.scala 43:21:@2833.4]
    .io_s(FA_24_io_s),
    .io_cout(FA_24_io_cout),
    .io_a(FA_24_io_a),
    .io_b(FA_24_io_b),
    .io_cin(FA_24_io_cin)
  );
  FA FA_25 ( // @[RA_Mul.scala 43:21:@2843.4]
    .io_s(FA_25_io_s),
    .io_cout(FA_25_io_cout),
    .io_a(FA_25_io_a),
    .io_b(FA_25_io_b),
    .io_cin(FA_25_io_cin)
  );
  FA FA_26 ( // @[RA_Mul.scala 43:21:@2853.4]
    .io_s(FA_26_io_s),
    .io_cout(FA_26_io_cout),
    .io_a(FA_26_io_a),
    .io_b(FA_26_io_b),
    .io_cin(FA_26_io_cin)
  );
  FA FA_27 ( // @[RA_Mul.scala 43:21:@2863.4]
    .io_s(FA_27_io_s),
    .io_cout(FA_27_io_cout),
    .io_a(FA_27_io_a),
    .io_b(FA_27_io_b),
    .io_cin(FA_27_io_cin)
  );
  FA FA_28 ( // @[RA_Mul.scala 43:21:@2880.4]
    .io_s(FA_28_io_s),
    .io_cout(FA_28_io_cout),
    .io_a(FA_28_io_a),
    .io_b(FA_28_io_b),
    .io_cin(FA_28_io_cin)
  );
  assign io_matrix_o_0_0 = io_matrix_i_0_0; // @[RA_Mul.scala 341:21:@2576.4]
  assign io_matrix_o_0_1 = HA_io_s; // @[RA_Mul.scala 22:7:@2585.4]
  assign io_matrix_o_0_2 = io_matrix_i_0_2; // @[RA_Mul.scala 347:21:@2590.4]
  assign io_matrix_o_0_3 = FA_io_s; // @[RA_Mul.scala 47:7:@2599.4]
  assign io_matrix_o_0_4 = io_matrix_i_0_4; // @[RA_Mul.scala 353:21:@2604.4]
  assign io_matrix_o_0_5 = io_matrix_i_0_5; // @[RA_Mul.scala 357:21:@2607.4]
  assign io_matrix_o_0_6 = FA_1_io_s; // @[RA_Mul.scala 47:7:@2617.4]
  assign io_matrix_o_0_7 = FA_2_io_s; // @[RA_Mul.scala 47:7:@2628.4]
  assign io_matrix_o_0_8 = FA_3_io_s; // @[RA_Mul.scala 47:7:@2638.4]
  assign io_matrix_o_0_9 = FA_4_io_s; // @[RA_Mul.scala 47:7:@2648.4]
  assign io_matrix_o_0_10 = FA_5_io_s; // @[RA_Mul.scala 47:7:@2658.4]
  assign io_matrix_o_0_11 = FA_6_io_s; // @[RA_Mul.scala 47:7:@2668.4]
  assign io_matrix_o_0_12 = FA_7_io_s; // @[RA_Mul.scala 47:7:@2678.4]
  assign io_matrix_o_0_13 = FA_9_io_s; // @[RA_Mul.scala 47:7:@2695.4]
  assign io_matrix_o_0_14 = FA_10_io_s; // @[RA_Mul.scala 47:7:@2710.4]
  assign io_matrix_o_0_15 = FA_11_io_s; // @[RA_Mul.scala 47:7:@2725.4]
  assign io_matrix_o_0_16 = FA_13_io_s; // @[RA_Mul.scala 47:7:@2741.4]
  assign io_matrix_o_0_17 = FA_15_io_s; // @[RA_Mul.scala 47:7:@2757.4]
  assign io_matrix_o_0_18 = FA_17_io_s; // @[RA_Mul.scala 47:7:@2773.4]
  assign io_matrix_o_0_19 = FA_19_io_s; // @[RA_Mul.scala 47:7:@2789.4]
  assign io_matrix_o_0_20 = FA_21_io_s; // @[RA_Mul.scala 47:7:@2805.4]
  assign io_matrix_o_0_21 = FA_22_io_s; // @[RA_Mul.scala 47:7:@2820.4]
  assign io_matrix_o_0_22 = FA_23_io_s; // @[RA_Mul.scala 47:7:@2829.4]
  assign io_matrix_o_0_23 = FA_24_io_s; // @[RA_Mul.scala 47:7:@2839.4]
  assign io_matrix_o_0_24 = FA_25_io_s; // @[RA_Mul.scala 47:7:@2849.4]
  assign io_matrix_o_0_25 = FA_26_io_s; // @[RA_Mul.scala 47:7:@2859.4]
  assign io_matrix_o_0_26 = FA_27_io_s; // @[RA_Mul.scala 47:7:@2869.4]
  assign io_matrix_o_0_27 = io_matrix_i_0_27; // @[RA_Mul.scala 422:22:@2873.4]
  assign io_matrix_o_0_28 = io_matrix_i_0_28; // @[RA_Mul.scala 426:22:@2876.4]
  assign io_matrix_o_0_29 = FA_28_io_s; // @[RA_Mul.scala 47:7:@2886.4]
  assign io_matrix_o_0_30 = io_matrix_i_0_30; // @[RA_Mul.scala 433:22:@2891.4]
  assign io_matrix_o_0_31 = io_matrix_i_0_31; // @[RA_Mul.scala 437:22:@2894.4]
  assign io_matrix_o_1_2 = HA_io_cout; // @[RA_Mul.scala 23:10:@2586.4]
  assign io_matrix_o_1_4 = FA_io_cout; // @[RA_Mul.scala 48:10:@2600.4]
  assign io_matrix_o_1_5 = io_matrix_i_1_5; // @[RA_Mul.scala 358:21:@2608.4]
  assign io_matrix_o_1_6 = io_matrix_i_3_6; // @[RA_Mul.scala 362:21:@2619.4]
  assign io_matrix_o_1_7 = FA_1_io_cout; // @[RA_Mul.scala 48:10:@2618.4]
  assign io_matrix_o_1_8 = FA_2_io_cout; // @[RA_Mul.scala 48:10:@2629.4]
  assign io_matrix_o_1_9 = FA_3_io_cout; // @[RA_Mul.scala 48:10:@2639.4]
  assign io_matrix_o_1_10 = FA_4_io_cout; // @[RA_Mul.scala 48:10:@2649.4]
  assign io_matrix_o_1_11 = FA_5_io_cout; // @[RA_Mul.scala 48:10:@2659.4]
  assign io_matrix_o_1_12 = FA_6_io_cout; // @[RA_Mul.scala 48:10:@2669.4]
  assign io_matrix_o_1_13 = FA_7_io_cout; // @[RA_Mul.scala 48:10:@2679.4]
  assign io_matrix_o_1_14 = FA_9_io_cout; // @[RA_Mul.scala 48:10:@2696.4]
  assign io_matrix_o_1_15 = FA_10_io_cout; // @[RA_Mul.scala 48:10:@2711.4]
  assign io_matrix_o_1_16 = FA_11_io_cout; // @[RA_Mul.scala 48:10:@2726.4]
  assign io_matrix_o_1_17 = FA_13_io_cout; // @[RA_Mul.scala 48:10:@2742.4]
  assign io_matrix_o_1_18 = FA_15_io_cout; // @[RA_Mul.scala 48:10:@2758.4]
  assign io_matrix_o_1_19 = FA_17_io_cout; // @[RA_Mul.scala 48:10:@2774.4]
  assign io_matrix_o_1_20 = FA_19_io_cout; // @[RA_Mul.scala 48:10:@2790.4]
  assign io_matrix_o_1_21 = FA_21_io_cout; // @[RA_Mul.scala 48:10:@2806.4]
  assign io_matrix_o_1_22 = FA_22_io_cout; // @[RA_Mul.scala 48:10:@2821.4]
  assign io_matrix_o_1_23 = FA_23_io_cout; // @[RA_Mul.scala 48:10:@2830.4]
  assign io_matrix_o_1_24 = FA_24_io_cout; // @[RA_Mul.scala 48:10:@2840.4]
  assign io_matrix_o_1_25 = FA_25_io_cout; // @[RA_Mul.scala 48:10:@2850.4]
  assign io_matrix_o_1_26 = FA_26_io_cout; // @[RA_Mul.scala 48:10:@2860.4]
  assign io_matrix_o_1_27 = FA_27_io_cout; // @[RA_Mul.scala 48:10:@2870.4]
  assign io_matrix_o_1_28 = io_matrix_i_1_28; // @[RA_Mul.scala 427:22:@2877.4]
  assign io_matrix_o_1_30 = FA_28_io_cout; // @[RA_Mul.scala 48:10:@2887.4]
  assign io_matrix_o_2_4 = io_matrix_i_1_4; // @[RA_Mul.scala 354:21:@2605.4]
  assign io_matrix_o_2_9 = io_matrix_i_3_9; // @[RA_Mul.scala 372:21:@2650.4]
  assign io_matrix_o_2_10 = io_matrix_i_3_10; // @[RA_Mul.scala 376:22:@2660.4]
  assign io_matrix_o_2_11 = io_matrix_i_3_11; // @[RA_Mul.scala 380:22:@2670.4]
  assign io_matrix_o_2_12 = FA_8_io_s; // @[RA_Mul.scala 47:7:@2686.4]
  assign io_matrix_o_2_13 = HA_1_io_s; // @[RA_Mul.scala 22:7:@2702.4]
  assign io_matrix_o_2_14 = HA_2_io_s; // @[RA_Mul.scala 22:7:@2717.4]
  assign io_matrix_o_2_15 = FA_12_io_s; // @[RA_Mul.scala 47:7:@2733.4]
  assign io_matrix_o_2_16 = FA_14_io_s; // @[RA_Mul.scala 47:7:@2749.4]
  assign io_matrix_o_2_17 = FA_16_io_s; // @[RA_Mul.scala 47:7:@2765.4]
  assign io_matrix_o_2_18 = FA_18_io_s; // @[RA_Mul.scala 47:7:@2781.4]
  assign io_matrix_o_2_19 = FA_20_io_s; // @[RA_Mul.scala 47:7:@2797.4]
  assign io_matrix_o_2_20 = HA_3_io_s; // @[RA_Mul.scala 22:7:@2812.4]
  assign io_matrix_o_2_21 = io_matrix_i_3_21; // @[RA_Mul.scala 402:22:@2822.4]
  assign io_matrix_o_2_22 = io_matrix_i_3_22; // @[RA_Mul.scala 405:22:@2831.4]
  assign io_matrix_o_2_23 = io_matrix_i_3_23; // @[RA_Mul.scala 409:22:@2841.4]
  assign io_matrix_o_2_24 = io_matrix_i_3_24; // @[RA_Mul.scala 413:22:@2851.4]
  assign io_matrix_o_2_27 = io_matrix_i_1_27; // @[RA_Mul.scala 423:22:@2874.4]
  assign io_matrix_o_2_30 = io_matrix_i_1_30; // @[RA_Mul.scala 434:22:@2892.4]
  assign io_matrix_o_3_9 = io_matrix_i_4_9; // @[RA_Mul.scala 373:21:@2651.4]
  assign io_matrix_o_3_13 = FA_8_io_cout; // @[RA_Mul.scala 48:10:@2687.4]
  assign io_matrix_o_3_14 = HA_1_io_cout; // @[RA_Mul.scala 23:10:@2703.4]
  assign io_matrix_o_3_15 = HA_2_io_cout; // @[RA_Mul.scala 23:10:@2718.4]
  assign io_matrix_o_3_16 = FA_12_io_cout; // @[RA_Mul.scala 48:10:@2734.4]
  assign io_matrix_o_3_17 = FA_14_io_cout; // @[RA_Mul.scala 48:10:@2750.4]
  assign io_matrix_o_3_18 = FA_16_io_cout; // @[RA_Mul.scala 48:10:@2766.4]
  assign io_matrix_o_3_19 = FA_18_io_cout; // @[RA_Mul.scala 48:10:@2782.4]
  assign io_matrix_o_3_20 = FA_20_io_cout; // @[RA_Mul.scala 48:10:@2798.4]
  assign io_matrix_o_3_21 = HA_3_io_cout; // @[RA_Mul.scala 23:10:@2813.4]
  assign io_matrix_o_3_23 = io_matrix_i_4_23; // @[RA_Mul.scala 410:22:@2842.4]
  assign HA_io_a = io_matrix_i_0_1; // @[RA_Mul.scala 20:14:@2583.4]
  assign HA_io_b = io_matrix_i_1_1; // @[RA_Mul.scala 21:14:@2584.4]
  assign FA_io_a = io_matrix_i_0_3; // @[RA_Mul.scala 44:14:@2596.4]
  assign FA_io_b = io_matrix_i_1_3; // @[RA_Mul.scala 45:14:@2597.4]
  assign FA_io_cin = io_matrix_i_2_3; // @[RA_Mul.scala 46:16:@2598.4]
  assign FA_1_io_a = io_matrix_i_0_6; // @[RA_Mul.scala 44:14:@2614.4]
  assign FA_1_io_b = io_matrix_i_1_6; // @[RA_Mul.scala 45:14:@2615.4]
  assign FA_1_io_cin = io_matrix_i_2_6; // @[RA_Mul.scala 46:16:@2616.4]
  assign FA_2_io_a = io_matrix_i_0_7; // @[RA_Mul.scala 44:14:@2625.4]
  assign FA_2_io_b = io_matrix_i_1_7; // @[RA_Mul.scala 45:14:@2626.4]
  assign FA_2_io_cin = io_matrix_i_2_7; // @[RA_Mul.scala 46:16:@2627.4]
  assign FA_3_io_a = io_matrix_i_0_8; // @[RA_Mul.scala 44:14:@2635.4]
  assign FA_3_io_b = io_matrix_i_1_8; // @[RA_Mul.scala 45:14:@2636.4]
  assign FA_3_io_cin = io_matrix_i_2_8; // @[RA_Mul.scala 46:16:@2637.4]
  assign FA_4_io_a = io_matrix_i_0_9; // @[RA_Mul.scala 44:14:@2645.4]
  assign FA_4_io_b = io_matrix_i_1_9; // @[RA_Mul.scala 45:14:@2646.4]
  assign FA_4_io_cin = io_matrix_i_2_9; // @[RA_Mul.scala 46:16:@2647.4]
  assign FA_5_io_a = io_matrix_i_0_10; // @[RA_Mul.scala 44:14:@2655.4]
  assign FA_5_io_b = io_matrix_i_1_10; // @[RA_Mul.scala 45:14:@2656.4]
  assign FA_5_io_cin = io_matrix_i_2_10; // @[RA_Mul.scala 46:16:@2657.4]
  assign FA_6_io_a = io_matrix_i_0_11; // @[RA_Mul.scala 44:14:@2665.4]
  assign FA_6_io_b = io_matrix_i_1_11; // @[RA_Mul.scala 45:14:@2666.4]
  assign FA_6_io_cin = io_matrix_i_2_11; // @[RA_Mul.scala 46:16:@2667.4]
  assign FA_7_io_a = io_matrix_i_0_12; // @[RA_Mul.scala 44:14:@2675.4]
  assign FA_7_io_b = io_matrix_i_1_12; // @[RA_Mul.scala 45:14:@2676.4]
  assign FA_7_io_cin = io_matrix_i_2_12; // @[RA_Mul.scala 46:16:@2677.4]
  assign FA_8_io_a = io_matrix_i_3_12; // @[RA_Mul.scala 44:14:@2683.4]
  assign FA_8_io_b = io_matrix_i_4_12; // @[RA_Mul.scala 45:14:@2684.4]
  assign FA_8_io_cin = io_matrix_i_5_12; // @[RA_Mul.scala 46:16:@2685.4]
  assign FA_9_io_a = io_matrix_i_0_13; // @[RA_Mul.scala 44:14:@2692.4]
  assign FA_9_io_b = io_matrix_i_1_13; // @[RA_Mul.scala 45:14:@2693.4]
  assign FA_9_io_cin = io_matrix_i_2_13; // @[RA_Mul.scala 46:16:@2694.4]
  assign HA_1_io_a = io_matrix_i_3_13; // @[RA_Mul.scala 20:14:@2700.4]
  assign HA_1_io_b = io_matrix_i_4_13; // @[RA_Mul.scala 21:14:@2701.4]
  assign FA_10_io_a = io_matrix_i_0_14; // @[RA_Mul.scala 44:14:@2707.4]
  assign FA_10_io_b = io_matrix_i_1_14; // @[RA_Mul.scala 45:14:@2708.4]
  assign FA_10_io_cin = io_matrix_i_2_14; // @[RA_Mul.scala 46:16:@2709.4]
  assign HA_2_io_a = io_matrix_i_3_14; // @[RA_Mul.scala 20:14:@2715.4]
  assign HA_2_io_b = io_matrix_i_4_14; // @[RA_Mul.scala 21:14:@2716.4]
  assign FA_11_io_a = io_matrix_i_0_15; // @[RA_Mul.scala 44:14:@2722.4]
  assign FA_11_io_b = io_matrix_i_1_15; // @[RA_Mul.scala 45:14:@2723.4]
  assign FA_11_io_cin = io_matrix_i_2_15; // @[RA_Mul.scala 46:16:@2724.4]
  assign FA_12_io_a = io_matrix_i_3_15; // @[RA_Mul.scala 44:14:@2730.4]
  assign FA_12_io_b = io_matrix_i_4_15; // @[RA_Mul.scala 45:14:@2731.4]
  assign FA_12_io_cin = io_matrix_i_5_15; // @[RA_Mul.scala 46:16:@2732.4]
  assign FA_13_io_a = io_matrix_i_0_16; // @[RA_Mul.scala 44:14:@2738.4]
  assign FA_13_io_b = io_matrix_i_1_16; // @[RA_Mul.scala 45:14:@2739.4]
  assign FA_13_io_cin = io_matrix_i_2_16; // @[RA_Mul.scala 46:16:@2740.4]
  assign FA_14_io_a = io_matrix_i_3_16; // @[RA_Mul.scala 44:14:@2746.4]
  assign FA_14_io_b = io_matrix_i_4_16; // @[RA_Mul.scala 45:14:@2747.4]
  assign FA_14_io_cin = io_matrix_i_5_16; // @[RA_Mul.scala 46:16:@2748.4]
  assign FA_15_io_a = io_matrix_i_0_17; // @[RA_Mul.scala 44:14:@2754.4]
  assign FA_15_io_b = io_matrix_i_1_17; // @[RA_Mul.scala 45:14:@2755.4]
  assign FA_15_io_cin = io_matrix_i_2_17; // @[RA_Mul.scala 46:16:@2756.4]
  assign FA_16_io_a = io_matrix_i_3_17; // @[RA_Mul.scala 44:14:@2762.4]
  assign FA_16_io_b = io_matrix_i_4_17; // @[RA_Mul.scala 45:14:@2763.4]
  assign FA_16_io_cin = io_matrix_i_5_17; // @[RA_Mul.scala 46:16:@2764.4]
  assign FA_17_io_a = io_matrix_i_0_18; // @[RA_Mul.scala 44:14:@2770.4]
  assign FA_17_io_b = io_matrix_i_1_18; // @[RA_Mul.scala 45:14:@2771.4]
  assign FA_17_io_cin = io_matrix_i_2_18; // @[RA_Mul.scala 46:16:@2772.4]
  assign FA_18_io_a = io_matrix_i_3_18; // @[RA_Mul.scala 44:14:@2778.4]
  assign FA_18_io_b = io_matrix_i_4_18; // @[RA_Mul.scala 45:14:@2779.4]
  assign FA_18_io_cin = io_matrix_i_5_18; // @[RA_Mul.scala 46:16:@2780.4]
  assign FA_19_io_a = io_matrix_i_0_19; // @[RA_Mul.scala 44:14:@2786.4]
  assign FA_19_io_b = io_matrix_i_1_19; // @[RA_Mul.scala 45:14:@2787.4]
  assign FA_19_io_cin = io_matrix_i_2_19; // @[RA_Mul.scala 46:16:@2788.4]
  assign FA_20_io_a = io_matrix_i_3_19; // @[RA_Mul.scala 44:14:@2794.4]
  assign FA_20_io_b = io_matrix_i_4_19; // @[RA_Mul.scala 45:14:@2795.4]
  assign FA_20_io_cin = io_matrix_i_5_19; // @[RA_Mul.scala 46:16:@2796.4]
  assign FA_21_io_a = io_matrix_i_0_20; // @[RA_Mul.scala 44:14:@2802.4]
  assign FA_21_io_b = io_matrix_i_1_20; // @[RA_Mul.scala 45:14:@2803.4]
  assign FA_21_io_cin = io_matrix_i_2_20; // @[RA_Mul.scala 46:16:@2804.4]
  assign HA_3_io_a = io_matrix_i_3_20; // @[RA_Mul.scala 20:14:@2810.4]
  assign HA_3_io_b = io_matrix_i_4_20; // @[RA_Mul.scala 21:14:@2811.4]
  assign FA_22_io_a = io_matrix_i_0_21; // @[RA_Mul.scala 44:14:@2817.4]
  assign FA_22_io_b = io_matrix_i_1_21; // @[RA_Mul.scala 45:14:@2818.4]
  assign FA_22_io_cin = io_matrix_i_2_21; // @[RA_Mul.scala 46:16:@2819.4]
  assign FA_23_io_a = io_matrix_i_0_22; // @[RA_Mul.scala 44:14:@2826.4]
  assign FA_23_io_b = io_matrix_i_1_22; // @[RA_Mul.scala 45:14:@2827.4]
  assign FA_23_io_cin = io_matrix_i_2_22; // @[RA_Mul.scala 46:16:@2828.4]
  assign FA_24_io_a = io_matrix_i_0_23; // @[RA_Mul.scala 44:14:@2836.4]
  assign FA_24_io_b = io_matrix_i_1_23; // @[RA_Mul.scala 45:14:@2837.4]
  assign FA_24_io_cin = io_matrix_i_2_23; // @[RA_Mul.scala 46:16:@2838.4]
  assign FA_25_io_a = io_matrix_i_0_24; // @[RA_Mul.scala 44:14:@2846.4]
  assign FA_25_io_b = io_matrix_i_1_24; // @[RA_Mul.scala 45:14:@2847.4]
  assign FA_25_io_cin = io_matrix_i_2_24; // @[RA_Mul.scala 46:16:@2848.4]
  assign FA_26_io_a = io_matrix_i_0_25; // @[RA_Mul.scala 44:14:@2856.4]
  assign FA_26_io_b = io_matrix_i_1_25; // @[RA_Mul.scala 45:14:@2857.4]
  assign FA_26_io_cin = io_matrix_i_2_25; // @[RA_Mul.scala 46:16:@2858.4]
  assign FA_27_io_a = io_matrix_i_0_26; // @[RA_Mul.scala 44:14:@2866.4]
  assign FA_27_io_b = io_matrix_i_1_26; // @[RA_Mul.scala 45:14:@2867.4]
  assign FA_27_io_cin = io_matrix_i_2_26; // @[RA_Mul.scala 46:16:@2868.4]
  assign FA_28_io_a = io_matrix_i_0_29; // @[RA_Mul.scala 44:14:@2883.4]
  assign FA_28_io_b = io_matrix_i_1_29; // @[RA_Mul.scala 45:14:@2884.4]
  assign FA_28_io_cin = io_matrix_i_2_29; // @[RA_Mul.scala 46:16:@2885.4]
endmodule
module Reduction_3( // @[:@3194.2]
  output  io_matrix_o_0_0, // @[:@3197.4]
  output  io_matrix_o_0_1, // @[:@3197.4]
  output  io_matrix_o_0_2, // @[:@3197.4]
  output  io_matrix_o_0_3, // @[:@3197.4]
  output  io_matrix_o_0_4, // @[:@3197.4]
  output  io_matrix_o_0_5, // @[:@3197.4]
  output  io_matrix_o_0_6, // @[:@3197.4]
  output  io_matrix_o_0_7, // @[:@3197.4]
  output  io_matrix_o_0_8, // @[:@3197.4]
  output  io_matrix_o_0_9, // @[:@3197.4]
  output  io_matrix_o_0_10, // @[:@3197.4]
  output  io_matrix_o_0_11, // @[:@3197.4]
  output  io_matrix_o_0_12, // @[:@3197.4]
  output  io_matrix_o_0_13, // @[:@3197.4]
  output  io_matrix_o_0_14, // @[:@3197.4]
  output  io_matrix_o_0_15, // @[:@3197.4]
  output  io_matrix_o_0_16, // @[:@3197.4]
  output  io_matrix_o_0_17, // @[:@3197.4]
  output  io_matrix_o_0_18, // @[:@3197.4]
  output  io_matrix_o_0_19, // @[:@3197.4]
  output  io_matrix_o_0_20, // @[:@3197.4]
  output  io_matrix_o_0_21, // @[:@3197.4]
  output  io_matrix_o_0_22, // @[:@3197.4]
  output  io_matrix_o_0_23, // @[:@3197.4]
  output  io_matrix_o_0_24, // @[:@3197.4]
  output  io_matrix_o_0_25, // @[:@3197.4]
  output  io_matrix_o_0_26, // @[:@3197.4]
  output  io_matrix_o_0_27, // @[:@3197.4]
  output  io_matrix_o_0_28, // @[:@3197.4]
  output  io_matrix_o_0_29, // @[:@3197.4]
  output  io_matrix_o_0_30, // @[:@3197.4]
  output  io_matrix_o_0_31, // @[:@3197.4]
  output  io_matrix_o_1_3, // @[:@3197.4]
  output  io_matrix_o_1_5, // @[:@3197.4]
  output  io_matrix_o_1_6, // @[:@3197.4]
  output  io_matrix_o_1_7, // @[:@3197.4]
  output  io_matrix_o_1_8, // @[:@3197.4]
  output  io_matrix_o_1_9, // @[:@3197.4]
  output  io_matrix_o_1_10, // @[:@3197.4]
  output  io_matrix_o_1_11, // @[:@3197.4]
  output  io_matrix_o_1_12, // @[:@3197.4]
  output  io_matrix_o_1_13, // @[:@3197.4]
  output  io_matrix_o_1_14, // @[:@3197.4]
  output  io_matrix_o_1_15, // @[:@3197.4]
  output  io_matrix_o_1_16, // @[:@3197.4]
  output  io_matrix_o_1_17, // @[:@3197.4]
  output  io_matrix_o_1_18, // @[:@3197.4]
  output  io_matrix_o_1_19, // @[:@3197.4]
  output  io_matrix_o_1_20, // @[:@3197.4]
  output  io_matrix_o_1_21, // @[:@3197.4]
  output  io_matrix_o_1_22, // @[:@3197.4]
  output  io_matrix_o_1_23, // @[:@3197.4]
  output  io_matrix_o_1_24, // @[:@3197.4]
  output  io_matrix_o_1_25, // @[:@3197.4]
  output  io_matrix_o_1_26, // @[:@3197.4]
  output  io_matrix_o_1_28, // @[:@3197.4]
  output  io_matrix_o_1_31, // @[:@3197.4]
  output  io_matrix_o_2_5, // @[:@3197.4]
  output  io_matrix_o_2_13, // @[:@3197.4]
  output  io_matrix_o_2_14, // @[:@3197.4]
  output  io_matrix_o_2_15, // @[:@3197.4]
  output  io_matrix_o_2_16, // @[:@3197.4]
  output  io_matrix_o_2_17, // @[:@3197.4]
  output  io_matrix_o_2_18, // @[:@3197.4]
  output  io_matrix_o_2_19, // @[:@3197.4]
  output  io_matrix_o_2_20, // @[:@3197.4]
  output  io_matrix_o_2_21, // @[:@3197.4]
  output  io_matrix_o_2_23, // @[:@3197.4]
  output  io_matrix_o_2_25, // @[:@3197.4]
  output  io_matrix_o_2_28, // @[:@3197.4]
  input   io_matrix_i_0_0, // @[:@3197.4]
  input   io_matrix_i_0_1, // @[:@3197.4]
  input   io_matrix_i_0_2, // @[:@3197.4]
  input   io_matrix_i_0_3, // @[:@3197.4]
  input   io_matrix_i_0_4, // @[:@3197.4]
  input   io_matrix_i_0_5, // @[:@3197.4]
  input   io_matrix_i_0_6, // @[:@3197.4]
  input   io_matrix_i_0_7, // @[:@3197.4]
  input   io_matrix_i_0_8, // @[:@3197.4]
  input   io_matrix_i_0_9, // @[:@3197.4]
  input   io_matrix_i_0_10, // @[:@3197.4]
  input   io_matrix_i_0_11, // @[:@3197.4]
  input   io_matrix_i_0_12, // @[:@3197.4]
  input   io_matrix_i_0_13, // @[:@3197.4]
  input   io_matrix_i_0_14, // @[:@3197.4]
  input   io_matrix_i_0_15, // @[:@3197.4]
  input   io_matrix_i_0_16, // @[:@3197.4]
  input   io_matrix_i_0_17, // @[:@3197.4]
  input   io_matrix_i_0_18, // @[:@3197.4]
  input   io_matrix_i_0_19, // @[:@3197.4]
  input   io_matrix_i_0_20, // @[:@3197.4]
  input   io_matrix_i_0_21, // @[:@3197.4]
  input   io_matrix_i_0_22, // @[:@3197.4]
  input   io_matrix_i_0_23, // @[:@3197.4]
  input   io_matrix_i_0_24, // @[:@3197.4]
  input   io_matrix_i_0_25, // @[:@3197.4]
  input   io_matrix_i_0_26, // @[:@3197.4]
  input   io_matrix_i_0_27, // @[:@3197.4]
  input   io_matrix_i_0_28, // @[:@3197.4]
  input   io_matrix_i_0_29, // @[:@3197.4]
  input   io_matrix_i_0_30, // @[:@3197.4]
  input   io_matrix_i_0_31, // @[:@3197.4]
  input   io_matrix_i_1_2, // @[:@3197.4]
  input   io_matrix_i_1_4, // @[:@3197.4]
  input   io_matrix_i_1_5, // @[:@3197.4]
  input   io_matrix_i_1_6, // @[:@3197.4]
  input   io_matrix_i_1_7, // @[:@3197.4]
  input   io_matrix_i_1_8, // @[:@3197.4]
  input   io_matrix_i_1_9, // @[:@3197.4]
  input   io_matrix_i_1_10, // @[:@3197.4]
  input   io_matrix_i_1_11, // @[:@3197.4]
  input   io_matrix_i_1_12, // @[:@3197.4]
  input   io_matrix_i_1_13, // @[:@3197.4]
  input   io_matrix_i_1_14, // @[:@3197.4]
  input   io_matrix_i_1_15, // @[:@3197.4]
  input   io_matrix_i_1_16, // @[:@3197.4]
  input   io_matrix_i_1_17, // @[:@3197.4]
  input   io_matrix_i_1_18, // @[:@3197.4]
  input   io_matrix_i_1_19, // @[:@3197.4]
  input   io_matrix_i_1_20, // @[:@3197.4]
  input   io_matrix_i_1_21, // @[:@3197.4]
  input   io_matrix_i_1_22, // @[:@3197.4]
  input   io_matrix_i_1_23, // @[:@3197.4]
  input   io_matrix_i_1_24, // @[:@3197.4]
  input   io_matrix_i_1_25, // @[:@3197.4]
  input   io_matrix_i_1_26, // @[:@3197.4]
  input   io_matrix_i_1_27, // @[:@3197.4]
  input   io_matrix_i_1_28, // @[:@3197.4]
  input   io_matrix_i_1_30, // @[:@3197.4]
  input   io_matrix_i_2_4, // @[:@3197.4]
  input   io_matrix_i_2_9, // @[:@3197.4]
  input   io_matrix_i_2_10, // @[:@3197.4]
  input   io_matrix_i_2_11, // @[:@3197.4]
  input   io_matrix_i_2_12, // @[:@3197.4]
  input   io_matrix_i_2_13, // @[:@3197.4]
  input   io_matrix_i_2_14, // @[:@3197.4]
  input   io_matrix_i_2_15, // @[:@3197.4]
  input   io_matrix_i_2_16, // @[:@3197.4]
  input   io_matrix_i_2_17, // @[:@3197.4]
  input   io_matrix_i_2_18, // @[:@3197.4]
  input   io_matrix_i_2_19, // @[:@3197.4]
  input   io_matrix_i_2_20, // @[:@3197.4]
  input   io_matrix_i_2_21, // @[:@3197.4]
  input   io_matrix_i_2_22, // @[:@3197.4]
  input   io_matrix_i_2_23, // @[:@3197.4]
  input   io_matrix_i_2_24, // @[:@3197.4]
  input   io_matrix_i_2_27, // @[:@3197.4]
  input   io_matrix_i_2_30, // @[:@3197.4]
  input   io_matrix_i_3_9, // @[:@3197.4]
  input   io_matrix_i_3_13, // @[:@3197.4]
  input   io_matrix_i_3_14, // @[:@3197.4]
  input   io_matrix_i_3_15, // @[:@3197.4]
  input   io_matrix_i_3_16, // @[:@3197.4]
  input   io_matrix_i_3_17, // @[:@3197.4]
  input   io_matrix_i_3_18, // @[:@3197.4]
  input   io_matrix_i_3_19, // @[:@3197.4]
  input   io_matrix_i_3_20, // @[:@3197.4]
  input   io_matrix_i_3_21, // @[:@3197.4]
  input   io_matrix_i_3_23 // @[:@3197.4]
);
  wire  HA_io_s; // @[RA_Mul.scala 19:21:@3205.4]
  wire  HA_io_cout; // @[RA_Mul.scala 19:21:@3205.4]
  wire  HA_io_a; // @[RA_Mul.scala 19:21:@3205.4]
  wire  HA_io_b; // @[RA_Mul.scala 19:21:@3205.4]
  wire  FA_io_s; // @[RA_Mul.scala 43:21:@3216.4]
  wire  FA_io_cout; // @[RA_Mul.scala 43:21:@3216.4]
  wire  FA_io_a; // @[RA_Mul.scala 43:21:@3216.4]
  wire  FA_io_b; // @[RA_Mul.scala 43:21:@3216.4]
  wire  FA_io_cin; // @[RA_Mul.scala 43:21:@3216.4]
  wire  FA_1_io_s; // @[RA_Mul.scala 43:21:@3237.4]
  wire  FA_1_io_cout; // @[RA_Mul.scala 43:21:@3237.4]
  wire  FA_1_io_a; // @[RA_Mul.scala 43:21:@3237.4]
  wire  FA_1_io_b; // @[RA_Mul.scala 43:21:@3237.4]
  wire  FA_1_io_cin; // @[RA_Mul.scala 43:21:@3237.4]
  wire  FA_2_io_s; // @[RA_Mul.scala 43:21:@3247.4]
  wire  FA_2_io_cout; // @[RA_Mul.scala 43:21:@3247.4]
  wire  FA_2_io_a; // @[RA_Mul.scala 43:21:@3247.4]
  wire  FA_2_io_b; // @[RA_Mul.scala 43:21:@3247.4]
  wire  FA_2_io_cin; // @[RA_Mul.scala 43:21:@3247.4]
  wire  FA_3_io_s; // @[RA_Mul.scala 43:21:@3256.4]
  wire  FA_3_io_cout; // @[RA_Mul.scala 43:21:@3256.4]
  wire  FA_3_io_a; // @[RA_Mul.scala 43:21:@3256.4]
  wire  FA_3_io_b; // @[RA_Mul.scala 43:21:@3256.4]
  wire  FA_3_io_cin; // @[RA_Mul.scala 43:21:@3256.4]
  wire  FA_4_io_s; // @[RA_Mul.scala 43:21:@3265.4]
  wire  FA_4_io_cout; // @[RA_Mul.scala 43:21:@3265.4]
  wire  FA_4_io_a; // @[RA_Mul.scala 43:21:@3265.4]
  wire  FA_4_io_b; // @[RA_Mul.scala 43:21:@3265.4]
  wire  FA_4_io_cin; // @[RA_Mul.scala 43:21:@3265.4]
  wire  FA_5_io_s; // @[RA_Mul.scala 43:21:@3274.4]
  wire  FA_5_io_cout; // @[RA_Mul.scala 43:21:@3274.4]
  wire  FA_5_io_a; // @[RA_Mul.scala 43:21:@3274.4]
  wire  FA_5_io_b; // @[RA_Mul.scala 43:21:@3274.4]
  wire  FA_5_io_cin; // @[RA_Mul.scala 43:21:@3274.4]
  wire  FA_6_io_s; // @[RA_Mul.scala 43:21:@3283.4]
  wire  FA_6_io_cout; // @[RA_Mul.scala 43:21:@3283.4]
  wire  FA_6_io_a; // @[RA_Mul.scala 43:21:@3283.4]
  wire  FA_6_io_b; // @[RA_Mul.scala 43:21:@3283.4]
  wire  FA_6_io_cin; // @[RA_Mul.scala 43:21:@3283.4]
  wire  FA_7_io_s; // @[RA_Mul.scala 43:21:@3292.4]
  wire  FA_7_io_cout; // @[RA_Mul.scala 43:21:@3292.4]
  wire  FA_7_io_a; // @[RA_Mul.scala 43:21:@3292.4]
  wire  FA_7_io_b; // @[RA_Mul.scala 43:21:@3292.4]
  wire  FA_7_io_cin; // @[RA_Mul.scala 43:21:@3292.4]
  wire  FA_8_io_s; // @[RA_Mul.scala 43:21:@3301.4]
  wire  FA_8_io_cout; // @[RA_Mul.scala 43:21:@3301.4]
  wire  FA_8_io_a; // @[RA_Mul.scala 43:21:@3301.4]
  wire  FA_8_io_b; // @[RA_Mul.scala 43:21:@3301.4]
  wire  FA_8_io_cin; // @[RA_Mul.scala 43:21:@3301.4]
  wire  FA_9_io_s; // @[RA_Mul.scala 43:21:@3310.4]
  wire  FA_9_io_cout; // @[RA_Mul.scala 43:21:@3310.4]
  wire  FA_9_io_a; // @[RA_Mul.scala 43:21:@3310.4]
  wire  FA_9_io_b; // @[RA_Mul.scala 43:21:@3310.4]
  wire  FA_9_io_cin; // @[RA_Mul.scala 43:21:@3310.4]
  wire  FA_10_io_s; // @[RA_Mul.scala 43:21:@3319.4]
  wire  FA_10_io_cout; // @[RA_Mul.scala 43:21:@3319.4]
  wire  FA_10_io_a; // @[RA_Mul.scala 43:21:@3319.4]
  wire  FA_10_io_b; // @[RA_Mul.scala 43:21:@3319.4]
  wire  FA_10_io_cin; // @[RA_Mul.scala 43:21:@3319.4]
  wire  FA_11_io_s; // @[RA_Mul.scala 43:21:@3328.4]
  wire  FA_11_io_cout; // @[RA_Mul.scala 43:21:@3328.4]
  wire  FA_11_io_a; // @[RA_Mul.scala 43:21:@3328.4]
  wire  FA_11_io_b; // @[RA_Mul.scala 43:21:@3328.4]
  wire  FA_11_io_cin; // @[RA_Mul.scala 43:21:@3328.4]
  wire  FA_12_io_s; // @[RA_Mul.scala 43:21:@3337.4]
  wire  FA_12_io_cout; // @[RA_Mul.scala 43:21:@3337.4]
  wire  FA_12_io_a; // @[RA_Mul.scala 43:21:@3337.4]
  wire  FA_12_io_b; // @[RA_Mul.scala 43:21:@3337.4]
  wire  FA_12_io_cin; // @[RA_Mul.scala 43:21:@3337.4]
  wire  FA_13_io_s; // @[RA_Mul.scala 43:21:@3346.4]
  wire  FA_13_io_cout; // @[RA_Mul.scala 43:21:@3346.4]
  wire  FA_13_io_a; // @[RA_Mul.scala 43:21:@3346.4]
  wire  FA_13_io_b; // @[RA_Mul.scala 43:21:@3346.4]
  wire  FA_13_io_cin; // @[RA_Mul.scala 43:21:@3346.4]
  wire  FA_14_io_s; // @[RA_Mul.scala 43:21:@3355.4]
  wire  FA_14_io_cout; // @[RA_Mul.scala 43:21:@3355.4]
  wire  FA_14_io_a; // @[RA_Mul.scala 43:21:@3355.4]
  wire  FA_14_io_b; // @[RA_Mul.scala 43:21:@3355.4]
  wire  FA_14_io_cin; // @[RA_Mul.scala 43:21:@3355.4]
  wire  FA_15_io_s; // @[RA_Mul.scala 43:21:@3364.4]
  wire  FA_15_io_cout; // @[RA_Mul.scala 43:21:@3364.4]
  wire  FA_15_io_a; // @[RA_Mul.scala 43:21:@3364.4]
  wire  FA_15_io_b; // @[RA_Mul.scala 43:21:@3364.4]
  wire  FA_15_io_cin; // @[RA_Mul.scala 43:21:@3364.4]
  wire  FA_16_io_s; // @[RA_Mul.scala 43:21:@3373.4]
  wire  FA_16_io_cout; // @[RA_Mul.scala 43:21:@3373.4]
  wire  FA_16_io_a; // @[RA_Mul.scala 43:21:@3373.4]
  wire  FA_16_io_b; // @[RA_Mul.scala 43:21:@3373.4]
  wire  FA_16_io_cin; // @[RA_Mul.scala 43:21:@3373.4]
  wire  FA_17_io_s; // @[RA_Mul.scala 43:21:@3387.4]
  wire  FA_17_io_cout; // @[RA_Mul.scala 43:21:@3387.4]
  wire  FA_17_io_a; // @[RA_Mul.scala 43:21:@3387.4]
  wire  FA_17_io_b; // @[RA_Mul.scala 43:21:@3387.4]
  wire  FA_17_io_cin; // @[RA_Mul.scala 43:21:@3387.4]
  wire  FA_18_io_s; // @[RA_Mul.scala 43:21:@3402.4]
  wire  FA_18_io_cout; // @[RA_Mul.scala 43:21:@3402.4]
  wire  FA_18_io_a; // @[RA_Mul.scala 43:21:@3402.4]
  wire  FA_18_io_b; // @[RA_Mul.scala 43:21:@3402.4]
  wire  FA_18_io_cin; // @[RA_Mul.scala 43:21:@3402.4]
  HA HA ( // @[RA_Mul.scala 19:21:@3205.4]
    .io_s(HA_io_s),
    .io_cout(HA_io_cout),
    .io_a(HA_io_a),
    .io_b(HA_io_b)
  );
  FA FA ( // @[RA_Mul.scala 43:21:@3216.4]
    .io_s(FA_io_s),
    .io_cout(FA_io_cout),
    .io_a(FA_io_a),
    .io_b(FA_io_b),
    .io_cin(FA_io_cin)
  );
  FA FA_1 ( // @[RA_Mul.scala 43:21:@3237.4]
    .io_s(FA_1_io_s),
    .io_cout(FA_1_io_cout),
    .io_a(FA_1_io_a),
    .io_b(FA_1_io_b),
    .io_cin(FA_1_io_cin)
  );
  FA FA_2 ( // @[RA_Mul.scala 43:21:@3247.4]
    .io_s(FA_2_io_s),
    .io_cout(FA_2_io_cout),
    .io_a(FA_2_io_a),
    .io_b(FA_2_io_b),
    .io_cin(FA_2_io_cin)
  );
  FA FA_3 ( // @[RA_Mul.scala 43:21:@3256.4]
    .io_s(FA_3_io_s),
    .io_cout(FA_3_io_cout),
    .io_a(FA_3_io_a),
    .io_b(FA_3_io_b),
    .io_cin(FA_3_io_cin)
  );
  FA FA_4 ( // @[RA_Mul.scala 43:21:@3265.4]
    .io_s(FA_4_io_s),
    .io_cout(FA_4_io_cout),
    .io_a(FA_4_io_a),
    .io_b(FA_4_io_b),
    .io_cin(FA_4_io_cin)
  );
  FA FA_5 ( // @[RA_Mul.scala 43:21:@3274.4]
    .io_s(FA_5_io_s),
    .io_cout(FA_5_io_cout),
    .io_a(FA_5_io_a),
    .io_b(FA_5_io_b),
    .io_cin(FA_5_io_cin)
  );
  FA FA_6 ( // @[RA_Mul.scala 43:21:@3283.4]
    .io_s(FA_6_io_s),
    .io_cout(FA_6_io_cout),
    .io_a(FA_6_io_a),
    .io_b(FA_6_io_b),
    .io_cin(FA_6_io_cin)
  );
  FA FA_7 ( // @[RA_Mul.scala 43:21:@3292.4]
    .io_s(FA_7_io_s),
    .io_cout(FA_7_io_cout),
    .io_a(FA_7_io_a),
    .io_b(FA_7_io_b),
    .io_cin(FA_7_io_cin)
  );
  FA FA_8 ( // @[RA_Mul.scala 43:21:@3301.4]
    .io_s(FA_8_io_s),
    .io_cout(FA_8_io_cout),
    .io_a(FA_8_io_a),
    .io_b(FA_8_io_b),
    .io_cin(FA_8_io_cin)
  );
  FA FA_9 ( // @[RA_Mul.scala 43:21:@3310.4]
    .io_s(FA_9_io_s),
    .io_cout(FA_9_io_cout),
    .io_a(FA_9_io_a),
    .io_b(FA_9_io_b),
    .io_cin(FA_9_io_cin)
  );
  FA FA_10 ( // @[RA_Mul.scala 43:21:@3319.4]
    .io_s(FA_10_io_s),
    .io_cout(FA_10_io_cout),
    .io_a(FA_10_io_a),
    .io_b(FA_10_io_b),
    .io_cin(FA_10_io_cin)
  );
  FA FA_11 ( // @[RA_Mul.scala 43:21:@3328.4]
    .io_s(FA_11_io_s),
    .io_cout(FA_11_io_cout),
    .io_a(FA_11_io_a),
    .io_b(FA_11_io_b),
    .io_cin(FA_11_io_cin)
  );
  FA FA_12 ( // @[RA_Mul.scala 43:21:@3337.4]
    .io_s(FA_12_io_s),
    .io_cout(FA_12_io_cout),
    .io_a(FA_12_io_a),
    .io_b(FA_12_io_b),
    .io_cin(FA_12_io_cin)
  );
  FA FA_13 ( // @[RA_Mul.scala 43:21:@3346.4]
    .io_s(FA_13_io_s),
    .io_cout(FA_13_io_cout),
    .io_a(FA_13_io_a),
    .io_b(FA_13_io_b),
    .io_cin(FA_13_io_cin)
  );
  FA FA_14 ( // @[RA_Mul.scala 43:21:@3355.4]
    .io_s(FA_14_io_s),
    .io_cout(FA_14_io_cout),
    .io_a(FA_14_io_a),
    .io_b(FA_14_io_b),
    .io_cin(FA_14_io_cin)
  );
  FA FA_15 ( // @[RA_Mul.scala 43:21:@3364.4]
    .io_s(FA_15_io_s),
    .io_cout(FA_15_io_cout),
    .io_a(FA_15_io_a),
    .io_b(FA_15_io_b),
    .io_cin(FA_15_io_cin)
  );
  FA FA_16 ( // @[RA_Mul.scala 43:21:@3373.4]
    .io_s(FA_16_io_s),
    .io_cout(FA_16_io_cout),
    .io_a(FA_16_io_a),
    .io_b(FA_16_io_b),
    .io_cin(FA_16_io_cin)
  );
  FA FA_17 ( // @[RA_Mul.scala 43:21:@3387.4]
    .io_s(FA_17_io_s),
    .io_cout(FA_17_io_cout),
    .io_a(FA_17_io_a),
    .io_b(FA_17_io_b),
    .io_cin(FA_17_io_cin)
  );
  FA FA_18 ( // @[RA_Mul.scala 43:21:@3402.4]
    .io_s(FA_18_io_s),
    .io_cout(FA_18_io_cout),
    .io_a(FA_18_io_a),
    .io_b(FA_18_io_b),
    .io_cin(FA_18_io_cin)
  );
  assign io_matrix_o_0_0 = io_matrix_i_0_0; // @[RA_Mul.scala 463:21:@3199.4]
  assign io_matrix_o_0_1 = io_matrix_i_0_1; // @[RA_Mul.scala 466:21:@3202.4]
  assign io_matrix_o_0_2 = HA_io_s; // @[RA_Mul.scala 22:7:@3210.4]
  assign io_matrix_o_0_3 = io_matrix_i_0_3; // @[RA_Mul.scala 472:21:@3214.4]
  assign io_matrix_o_0_4 = FA_io_s; // @[RA_Mul.scala 47:7:@3222.4]
  assign io_matrix_o_0_5 = io_matrix_i_0_5; // @[RA_Mul.scala 478:21:@3226.4]
  assign io_matrix_o_0_6 = io_matrix_i_0_6; // @[RA_Mul.scala 482:23:@3228.4]
  assign io_matrix_o_0_7 = io_matrix_i_0_7; // @[RA_Mul.scala 482:23:@3231.4]
  assign io_matrix_o_0_8 = io_matrix_i_0_8; // @[RA_Mul.scala 482:23:@3234.4]
  assign io_matrix_o_0_9 = FA_1_io_s; // @[RA_Mul.scala 47:7:@3243.4]
  assign io_matrix_o_0_10 = FA_2_io_s; // @[RA_Mul.scala 47:7:@3253.4]
  assign io_matrix_o_0_11 = FA_3_io_s; // @[RA_Mul.scala 47:7:@3262.4]
  assign io_matrix_o_0_12 = FA_4_io_s; // @[RA_Mul.scala 47:7:@3271.4]
  assign io_matrix_o_0_13 = FA_5_io_s; // @[RA_Mul.scala 47:7:@3280.4]
  assign io_matrix_o_0_14 = FA_6_io_s; // @[RA_Mul.scala 47:7:@3289.4]
  assign io_matrix_o_0_15 = FA_7_io_s; // @[RA_Mul.scala 47:7:@3298.4]
  assign io_matrix_o_0_16 = FA_8_io_s; // @[RA_Mul.scala 47:7:@3307.4]
  assign io_matrix_o_0_17 = FA_9_io_s; // @[RA_Mul.scala 47:7:@3316.4]
  assign io_matrix_o_0_18 = FA_10_io_s; // @[RA_Mul.scala 47:7:@3325.4]
  assign io_matrix_o_0_19 = FA_11_io_s; // @[RA_Mul.scala 47:7:@3334.4]
  assign io_matrix_o_0_20 = FA_12_io_s; // @[RA_Mul.scala 47:7:@3343.4]
  assign io_matrix_o_0_21 = FA_13_io_s; // @[RA_Mul.scala 47:7:@3352.4]
  assign io_matrix_o_0_22 = FA_14_io_s; // @[RA_Mul.scala 47:7:@3361.4]
  assign io_matrix_o_0_23 = FA_15_io_s; // @[RA_Mul.scala 47:7:@3370.4]
  assign io_matrix_o_0_24 = FA_16_io_s; // @[RA_Mul.scala 47:7:@3379.4]
  assign io_matrix_o_0_25 = io_matrix_i_0_25; // @[RA_Mul.scala 510:22:@3382.4]
  assign io_matrix_o_0_26 = io_matrix_i_0_26; // @[RA_Mul.scala 513:22:@3384.4]
  assign io_matrix_o_0_27 = FA_17_io_s; // @[RA_Mul.scala 47:7:@3393.4]
  assign io_matrix_o_0_28 = io_matrix_i_0_28; // @[RA_Mul.scala 520:22:@3397.4]
  assign io_matrix_o_0_29 = io_matrix_i_0_29; // @[RA_Mul.scala 523:22:@3399.4]
  assign io_matrix_o_0_30 = FA_18_io_s; // @[RA_Mul.scala 47:7:@3408.4]
  assign io_matrix_o_0_31 = io_matrix_i_0_31; // @[RA_Mul.scala 529:22:@3412.4]
  assign io_matrix_o_1_3 = HA_io_cout; // @[RA_Mul.scala 23:10:@3211.4]
  assign io_matrix_o_1_5 = FA_io_cout; // @[RA_Mul.scala 48:10:@3223.4]
  assign io_matrix_o_1_6 = io_matrix_i_1_6; // @[RA_Mul.scala 483:23:@3229.4]
  assign io_matrix_o_1_7 = io_matrix_i_1_7; // @[RA_Mul.scala 483:23:@3232.4]
  assign io_matrix_o_1_8 = io_matrix_i_1_8; // @[RA_Mul.scala 483:23:@3235.4]
  assign io_matrix_o_1_9 = io_matrix_i_3_9; // @[RA_Mul.scala 488:21:@3245.4]
  assign io_matrix_o_1_10 = FA_1_io_cout; // @[RA_Mul.scala 48:10:@3244.4]
  assign io_matrix_o_1_11 = FA_2_io_cout; // @[RA_Mul.scala 48:10:@3254.4]
  assign io_matrix_o_1_12 = FA_3_io_cout; // @[RA_Mul.scala 48:10:@3263.4]
  assign io_matrix_o_1_13 = FA_4_io_cout; // @[RA_Mul.scala 48:10:@3272.4]
  assign io_matrix_o_1_14 = FA_5_io_cout; // @[RA_Mul.scala 48:10:@3281.4]
  assign io_matrix_o_1_15 = FA_6_io_cout; // @[RA_Mul.scala 48:10:@3290.4]
  assign io_matrix_o_1_16 = FA_7_io_cout; // @[RA_Mul.scala 48:10:@3299.4]
  assign io_matrix_o_1_17 = FA_8_io_cout; // @[RA_Mul.scala 48:10:@3308.4]
  assign io_matrix_o_1_18 = FA_9_io_cout; // @[RA_Mul.scala 48:10:@3317.4]
  assign io_matrix_o_1_19 = FA_10_io_cout; // @[RA_Mul.scala 48:10:@3326.4]
  assign io_matrix_o_1_20 = FA_11_io_cout; // @[RA_Mul.scala 48:10:@3335.4]
  assign io_matrix_o_1_21 = FA_12_io_cout; // @[RA_Mul.scala 48:10:@3344.4]
  assign io_matrix_o_1_22 = FA_13_io_cout; // @[RA_Mul.scala 48:10:@3353.4]
  assign io_matrix_o_1_23 = FA_14_io_cout; // @[RA_Mul.scala 48:10:@3362.4]
  assign io_matrix_o_1_24 = FA_15_io_cout; // @[RA_Mul.scala 48:10:@3371.4]
  assign io_matrix_o_1_25 = FA_16_io_cout; // @[RA_Mul.scala 48:10:@3380.4]
  assign io_matrix_o_1_26 = io_matrix_i_1_26; // @[RA_Mul.scala 514:22:@3385.4]
  assign io_matrix_o_1_28 = FA_17_io_cout; // @[RA_Mul.scala 48:10:@3394.4]
  assign io_matrix_o_1_31 = FA_18_io_cout; // @[RA_Mul.scala 48:10:@3409.4]
  assign io_matrix_o_2_5 = io_matrix_i_1_5; // @[RA_Mul.scala 479:21:@3227.4]
  assign io_matrix_o_2_13 = io_matrix_i_3_13; // @[RA_Mul.scala 498:23:@3282.4]
  assign io_matrix_o_2_14 = io_matrix_i_3_14; // @[RA_Mul.scala 498:23:@3291.4]
  assign io_matrix_o_2_15 = io_matrix_i_3_15; // @[RA_Mul.scala 498:23:@3300.4]
  assign io_matrix_o_2_16 = io_matrix_i_3_16; // @[RA_Mul.scala 498:23:@3309.4]
  assign io_matrix_o_2_17 = io_matrix_i_3_17; // @[RA_Mul.scala 498:23:@3318.4]
  assign io_matrix_o_2_18 = io_matrix_i_3_18; // @[RA_Mul.scala 498:23:@3327.4]
  assign io_matrix_o_2_19 = io_matrix_i_3_19; // @[RA_Mul.scala 498:23:@3336.4]
  assign io_matrix_o_2_20 = io_matrix_i_3_20; // @[RA_Mul.scala 498:23:@3345.4]
  assign io_matrix_o_2_21 = io_matrix_i_3_21; // @[RA_Mul.scala 498:23:@3354.4]
  assign io_matrix_o_2_23 = io_matrix_i_3_23; // @[RA_Mul.scala 505:22:@3372.4]
  assign io_matrix_o_2_25 = io_matrix_i_1_25; // @[RA_Mul.scala 511:22:@3383.4]
  assign io_matrix_o_2_28 = io_matrix_i_1_28; // @[RA_Mul.scala 521:22:@3398.4]
  assign HA_io_a = io_matrix_i_0_2; // @[RA_Mul.scala 20:14:@3208.4]
  assign HA_io_b = io_matrix_i_1_2; // @[RA_Mul.scala 21:14:@3209.4]
  assign FA_io_a = io_matrix_i_0_4; // @[RA_Mul.scala 44:14:@3219.4]
  assign FA_io_b = io_matrix_i_1_4; // @[RA_Mul.scala 45:14:@3220.4]
  assign FA_io_cin = io_matrix_i_2_4; // @[RA_Mul.scala 46:16:@3221.4]
  assign FA_1_io_a = io_matrix_i_0_9; // @[RA_Mul.scala 44:14:@3240.4]
  assign FA_1_io_b = io_matrix_i_1_9; // @[RA_Mul.scala 45:14:@3241.4]
  assign FA_1_io_cin = io_matrix_i_2_9; // @[RA_Mul.scala 46:16:@3242.4]
  assign FA_2_io_a = io_matrix_i_0_10; // @[RA_Mul.scala 44:14:@3250.4]
  assign FA_2_io_b = io_matrix_i_1_10; // @[RA_Mul.scala 45:14:@3251.4]
  assign FA_2_io_cin = io_matrix_i_2_10; // @[RA_Mul.scala 46:16:@3252.4]
  assign FA_3_io_a = io_matrix_i_0_11; // @[RA_Mul.scala 44:14:@3259.4]
  assign FA_3_io_b = io_matrix_i_1_11; // @[RA_Mul.scala 45:14:@3260.4]
  assign FA_3_io_cin = io_matrix_i_2_11; // @[RA_Mul.scala 46:16:@3261.4]
  assign FA_4_io_a = io_matrix_i_0_12; // @[RA_Mul.scala 44:14:@3268.4]
  assign FA_4_io_b = io_matrix_i_1_12; // @[RA_Mul.scala 45:14:@3269.4]
  assign FA_4_io_cin = io_matrix_i_2_12; // @[RA_Mul.scala 46:16:@3270.4]
  assign FA_5_io_a = io_matrix_i_0_13; // @[RA_Mul.scala 44:14:@3277.4]
  assign FA_5_io_b = io_matrix_i_1_13; // @[RA_Mul.scala 45:14:@3278.4]
  assign FA_5_io_cin = io_matrix_i_2_13; // @[RA_Mul.scala 46:16:@3279.4]
  assign FA_6_io_a = io_matrix_i_0_14; // @[RA_Mul.scala 44:14:@3286.4]
  assign FA_6_io_b = io_matrix_i_1_14; // @[RA_Mul.scala 45:14:@3287.4]
  assign FA_6_io_cin = io_matrix_i_2_14; // @[RA_Mul.scala 46:16:@3288.4]
  assign FA_7_io_a = io_matrix_i_0_15; // @[RA_Mul.scala 44:14:@3295.4]
  assign FA_7_io_b = io_matrix_i_1_15; // @[RA_Mul.scala 45:14:@3296.4]
  assign FA_7_io_cin = io_matrix_i_2_15; // @[RA_Mul.scala 46:16:@3297.4]
  assign FA_8_io_a = io_matrix_i_0_16; // @[RA_Mul.scala 44:14:@3304.4]
  assign FA_8_io_b = io_matrix_i_1_16; // @[RA_Mul.scala 45:14:@3305.4]
  assign FA_8_io_cin = io_matrix_i_2_16; // @[RA_Mul.scala 46:16:@3306.4]
  assign FA_9_io_a = io_matrix_i_0_17; // @[RA_Mul.scala 44:14:@3313.4]
  assign FA_9_io_b = io_matrix_i_1_17; // @[RA_Mul.scala 45:14:@3314.4]
  assign FA_9_io_cin = io_matrix_i_2_17; // @[RA_Mul.scala 46:16:@3315.4]
  assign FA_10_io_a = io_matrix_i_0_18; // @[RA_Mul.scala 44:14:@3322.4]
  assign FA_10_io_b = io_matrix_i_1_18; // @[RA_Mul.scala 45:14:@3323.4]
  assign FA_10_io_cin = io_matrix_i_2_18; // @[RA_Mul.scala 46:16:@3324.4]
  assign FA_11_io_a = io_matrix_i_0_19; // @[RA_Mul.scala 44:14:@3331.4]
  assign FA_11_io_b = io_matrix_i_1_19; // @[RA_Mul.scala 45:14:@3332.4]
  assign FA_11_io_cin = io_matrix_i_2_19; // @[RA_Mul.scala 46:16:@3333.4]
  assign FA_12_io_a = io_matrix_i_0_20; // @[RA_Mul.scala 44:14:@3340.4]
  assign FA_12_io_b = io_matrix_i_1_20; // @[RA_Mul.scala 45:14:@3341.4]
  assign FA_12_io_cin = io_matrix_i_2_20; // @[RA_Mul.scala 46:16:@3342.4]
  assign FA_13_io_a = io_matrix_i_0_21; // @[RA_Mul.scala 44:14:@3349.4]
  assign FA_13_io_b = io_matrix_i_1_21; // @[RA_Mul.scala 45:14:@3350.4]
  assign FA_13_io_cin = io_matrix_i_2_21; // @[RA_Mul.scala 46:16:@3351.4]
  assign FA_14_io_a = io_matrix_i_0_22; // @[RA_Mul.scala 44:14:@3358.4]
  assign FA_14_io_b = io_matrix_i_1_22; // @[RA_Mul.scala 45:14:@3359.4]
  assign FA_14_io_cin = io_matrix_i_2_22; // @[RA_Mul.scala 46:16:@3360.4]
  assign FA_15_io_a = io_matrix_i_0_23; // @[RA_Mul.scala 44:14:@3367.4]
  assign FA_15_io_b = io_matrix_i_1_23; // @[RA_Mul.scala 45:14:@3368.4]
  assign FA_15_io_cin = io_matrix_i_2_23; // @[RA_Mul.scala 46:16:@3369.4]
  assign FA_16_io_a = io_matrix_i_0_24; // @[RA_Mul.scala 44:14:@3376.4]
  assign FA_16_io_b = io_matrix_i_1_24; // @[RA_Mul.scala 45:14:@3377.4]
  assign FA_16_io_cin = io_matrix_i_2_24; // @[RA_Mul.scala 46:16:@3378.4]
  assign FA_17_io_a = io_matrix_i_0_27; // @[RA_Mul.scala 44:14:@3390.4]
  assign FA_17_io_b = io_matrix_i_1_27; // @[RA_Mul.scala 45:14:@3391.4]
  assign FA_17_io_cin = io_matrix_i_2_27; // @[RA_Mul.scala 46:16:@3392.4]
  assign FA_18_io_a = io_matrix_i_0_30; // @[RA_Mul.scala 44:14:@3405.4]
  assign FA_18_io_b = io_matrix_i_1_30; // @[RA_Mul.scala 45:14:@3406.4]
  assign FA_18_io_cin = io_matrix_i_2_30; // @[RA_Mul.scala 46:16:@3407.4]
endmodule
module Reduction_4( // @[:@3720.2]
  output  io_matrix_o_0_0, // @[:@3723.4]
  output  io_matrix_o_0_1, // @[:@3723.4]
  output  io_matrix_o_0_2, // @[:@3723.4]
  output  io_matrix_o_0_3, // @[:@3723.4]
  output  io_matrix_o_0_4, // @[:@3723.4]
  output  io_matrix_o_0_5, // @[:@3723.4]
  output  io_matrix_o_0_6, // @[:@3723.4]
  output  io_matrix_o_0_7, // @[:@3723.4]
  output  io_matrix_o_0_8, // @[:@3723.4]
  output  io_matrix_o_0_9, // @[:@3723.4]
  output  io_matrix_o_0_10, // @[:@3723.4]
  output  io_matrix_o_0_11, // @[:@3723.4]
  output  io_matrix_o_0_12, // @[:@3723.4]
  output  io_matrix_o_0_13, // @[:@3723.4]
  output  io_matrix_o_0_14, // @[:@3723.4]
  output  io_matrix_o_0_15, // @[:@3723.4]
  output  io_matrix_o_0_16, // @[:@3723.4]
  output  io_matrix_o_0_17, // @[:@3723.4]
  output  io_matrix_o_0_18, // @[:@3723.4]
  output  io_matrix_o_0_19, // @[:@3723.4]
  output  io_matrix_o_0_20, // @[:@3723.4]
  output  io_matrix_o_0_21, // @[:@3723.4]
  output  io_matrix_o_0_22, // @[:@3723.4]
  output  io_matrix_o_0_23, // @[:@3723.4]
  output  io_matrix_o_0_24, // @[:@3723.4]
  output  io_matrix_o_0_25, // @[:@3723.4]
  output  io_matrix_o_0_26, // @[:@3723.4]
  output  io_matrix_o_0_27, // @[:@3723.4]
  output  io_matrix_o_0_28, // @[:@3723.4]
  output  io_matrix_o_0_29, // @[:@3723.4]
  output  io_matrix_o_0_30, // @[:@3723.4]
  output  io_matrix_o_0_31, // @[:@3723.4]
  output  io_matrix_o_1_4, // @[:@3723.4]
  output  io_matrix_o_1_6, // @[:@3723.4]
  output  io_matrix_o_1_7, // @[:@3723.4]
  output  io_matrix_o_1_8, // @[:@3723.4]
  output  io_matrix_o_1_9, // @[:@3723.4]
  output  io_matrix_o_1_10, // @[:@3723.4]
  output  io_matrix_o_1_11, // @[:@3723.4]
  output  io_matrix_o_1_12, // @[:@3723.4]
  output  io_matrix_o_1_13, // @[:@3723.4]
  output  io_matrix_o_1_14, // @[:@3723.4]
  output  io_matrix_o_1_15, // @[:@3723.4]
  output  io_matrix_o_1_16, // @[:@3723.4]
  output  io_matrix_o_1_17, // @[:@3723.4]
  output  io_matrix_o_1_18, // @[:@3723.4]
  output  io_matrix_o_1_19, // @[:@3723.4]
  output  io_matrix_o_1_20, // @[:@3723.4]
  output  io_matrix_o_1_21, // @[:@3723.4]
  output  io_matrix_o_1_22, // @[:@3723.4]
  output  io_matrix_o_1_23, // @[:@3723.4]
  output  io_matrix_o_1_24, // @[:@3723.4]
  output  io_matrix_o_1_25, // @[:@3723.4]
  output  io_matrix_o_1_26, // @[:@3723.4]
  output  io_matrix_o_1_27, // @[:@3723.4]
  output  io_matrix_o_1_29, // @[:@3723.4]
  output  io_matrix_o_1_31, // @[:@3723.4]
  input   io_matrix_i_0_0, // @[:@3723.4]
  input   io_matrix_i_0_1, // @[:@3723.4]
  input   io_matrix_i_0_2, // @[:@3723.4]
  input   io_matrix_i_0_3, // @[:@3723.4]
  input   io_matrix_i_0_4, // @[:@3723.4]
  input   io_matrix_i_0_5, // @[:@3723.4]
  input   io_matrix_i_0_6, // @[:@3723.4]
  input   io_matrix_i_0_7, // @[:@3723.4]
  input   io_matrix_i_0_8, // @[:@3723.4]
  input   io_matrix_i_0_9, // @[:@3723.4]
  input   io_matrix_i_0_10, // @[:@3723.4]
  input   io_matrix_i_0_11, // @[:@3723.4]
  input   io_matrix_i_0_12, // @[:@3723.4]
  input   io_matrix_i_0_13, // @[:@3723.4]
  input   io_matrix_i_0_14, // @[:@3723.4]
  input   io_matrix_i_0_15, // @[:@3723.4]
  input   io_matrix_i_0_16, // @[:@3723.4]
  input   io_matrix_i_0_17, // @[:@3723.4]
  input   io_matrix_i_0_18, // @[:@3723.4]
  input   io_matrix_i_0_19, // @[:@3723.4]
  input   io_matrix_i_0_20, // @[:@3723.4]
  input   io_matrix_i_0_21, // @[:@3723.4]
  input   io_matrix_i_0_22, // @[:@3723.4]
  input   io_matrix_i_0_23, // @[:@3723.4]
  input   io_matrix_i_0_24, // @[:@3723.4]
  input   io_matrix_i_0_25, // @[:@3723.4]
  input   io_matrix_i_0_26, // @[:@3723.4]
  input   io_matrix_i_0_27, // @[:@3723.4]
  input   io_matrix_i_0_28, // @[:@3723.4]
  input   io_matrix_i_0_29, // @[:@3723.4]
  input   io_matrix_i_0_30, // @[:@3723.4]
  input   io_matrix_i_0_31, // @[:@3723.4]
  input   io_matrix_i_1_3, // @[:@3723.4]
  input   io_matrix_i_1_5, // @[:@3723.4]
  input   io_matrix_i_1_6, // @[:@3723.4]
  input   io_matrix_i_1_7, // @[:@3723.4]
  input   io_matrix_i_1_8, // @[:@3723.4]
  input   io_matrix_i_1_9, // @[:@3723.4]
  input   io_matrix_i_1_10, // @[:@3723.4]
  input   io_matrix_i_1_11, // @[:@3723.4]
  input   io_matrix_i_1_12, // @[:@3723.4]
  input   io_matrix_i_1_13, // @[:@3723.4]
  input   io_matrix_i_1_14, // @[:@3723.4]
  input   io_matrix_i_1_15, // @[:@3723.4]
  input   io_matrix_i_1_16, // @[:@3723.4]
  input   io_matrix_i_1_17, // @[:@3723.4]
  input   io_matrix_i_1_18, // @[:@3723.4]
  input   io_matrix_i_1_19, // @[:@3723.4]
  input   io_matrix_i_1_20, // @[:@3723.4]
  input   io_matrix_i_1_21, // @[:@3723.4]
  input   io_matrix_i_1_22, // @[:@3723.4]
  input   io_matrix_i_1_23, // @[:@3723.4]
  input   io_matrix_i_1_24, // @[:@3723.4]
  input   io_matrix_i_1_25, // @[:@3723.4]
  input   io_matrix_i_1_26, // @[:@3723.4]
  input   io_matrix_i_1_28, // @[:@3723.4]
  input   io_matrix_i_1_31, // @[:@3723.4]
  input   io_matrix_i_2_5, // @[:@3723.4]
  input   io_matrix_i_2_13, // @[:@3723.4]
  input   io_matrix_i_2_14, // @[:@3723.4]
  input   io_matrix_i_2_15, // @[:@3723.4]
  input   io_matrix_i_2_16, // @[:@3723.4]
  input   io_matrix_i_2_17, // @[:@3723.4]
  input   io_matrix_i_2_18, // @[:@3723.4]
  input   io_matrix_i_2_19, // @[:@3723.4]
  input   io_matrix_i_2_20, // @[:@3723.4]
  input   io_matrix_i_2_21, // @[:@3723.4]
  input   io_matrix_i_2_23, // @[:@3723.4]
  input   io_matrix_i_2_25, // @[:@3723.4]
  input   io_matrix_i_2_28 // @[:@3723.4]
);
  wire  HA_io_s; // @[RA_Mul.scala 19:21:@3731.4]
  wire  HA_io_cout; // @[RA_Mul.scala 19:21:@3731.4]
  wire  HA_io_a; // @[RA_Mul.scala 19:21:@3731.4]
  wire  HA_io_b; // @[RA_Mul.scala 19:21:@3731.4]
  wire  FA_io_s; // @[RA_Mul.scala 43:21:@3740.4]
  wire  FA_io_cout; // @[RA_Mul.scala 43:21:@3740.4]
  wire  FA_io_a; // @[RA_Mul.scala 43:21:@3740.4]
  wire  FA_io_b; // @[RA_Mul.scala 43:21:@3740.4]
  wire  FA_io_cin; // @[RA_Mul.scala 43:21:@3740.4]
  wire  HA_1_io_s; // @[RA_Mul.scala 19:21:@3749.4]
  wire  HA_1_io_cout; // @[RA_Mul.scala 19:21:@3749.4]
  wire  HA_1_io_a; // @[RA_Mul.scala 19:21:@3749.4]
  wire  HA_1_io_b; // @[RA_Mul.scala 19:21:@3749.4]
  wire  HA_2_io_s; // @[RA_Mul.scala 19:21:@3756.4]
  wire  HA_2_io_cout; // @[RA_Mul.scala 19:21:@3756.4]
  wire  HA_2_io_a; // @[RA_Mul.scala 19:21:@3756.4]
  wire  HA_2_io_b; // @[RA_Mul.scala 19:21:@3756.4]
  wire  HA_3_io_s; // @[RA_Mul.scala 19:21:@3763.4]
  wire  HA_3_io_cout; // @[RA_Mul.scala 19:21:@3763.4]
  wire  HA_3_io_a; // @[RA_Mul.scala 19:21:@3763.4]
  wire  HA_3_io_b; // @[RA_Mul.scala 19:21:@3763.4]
  wire  HA_4_io_s; // @[RA_Mul.scala 19:21:@3770.4]
  wire  HA_4_io_cout; // @[RA_Mul.scala 19:21:@3770.4]
  wire  HA_4_io_a; // @[RA_Mul.scala 19:21:@3770.4]
  wire  HA_4_io_b; // @[RA_Mul.scala 19:21:@3770.4]
  wire  HA_5_io_s; // @[RA_Mul.scala 19:21:@3777.4]
  wire  HA_5_io_cout; // @[RA_Mul.scala 19:21:@3777.4]
  wire  HA_5_io_a; // @[RA_Mul.scala 19:21:@3777.4]
  wire  HA_5_io_b; // @[RA_Mul.scala 19:21:@3777.4]
  wire  HA_6_io_s; // @[RA_Mul.scala 19:21:@3784.4]
  wire  HA_6_io_cout; // @[RA_Mul.scala 19:21:@3784.4]
  wire  HA_6_io_a; // @[RA_Mul.scala 19:21:@3784.4]
  wire  HA_6_io_b; // @[RA_Mul.scala 19:21:@3784.4]
  wire  HA_7_io_s; // @[RA_Mul.scala 19:21:@3791.4]
  wire  HA_7_io_cout; // @[RA_Mul.scala 19:21:@3791.4]
  wire  HA_7_io_a; // @[RA_Mul.scala 19:21:@3791.4]
  wire  HA_7_io_b; // @[RA_Mul.scala 19:21:@3791.4]
  wire  FA_1_io_s; // @[RA_Mul.scala 43:21:@3798.4]
  wire  FA_1_io_cout; // @[RA_Mul.scala 43:21:@3798.4]
  wire  FA_1_io_a; // @[RA_Mul.scala 43:21:@3798.4]
  wire  FA_1_io_b; // @[RA_Mul.scala 43:21:@3798.4]
  wire  FA_1_io_cin; // @[RA_Mul.scala 43:21:@3798.4]
  wire  FA_2_io_s; // @[RA_Mul.scala 43:21:@3806.4]
  wire  FA_2_io_cout; // @[RA_Mul.scala 43:21:@3806.4]
  wire  FA_2_io_a; // @[RA_Mul.scala 43:21:@3806.4]
  wire  FA_2_io_b; // @[RA_Mul.scala 43:21:@3806.4]
  wire  FA_2_io_cin; // @[RA_Mul.scala 43:21:@3806.4]
  wire  FA_3_io_s; // @[RA_Mul.scala 43:21:@3814.4]
  wire  FA_3_io_cout; // @[RA_Mul.scala 43:21:@3814.4]
  wire  FA_3_io_a; // @[RA_Mul.scala 43:21:@3814.4]
  wire  FA_3_io_b; // @[RA_Mul.scala 43:21:@3814.4]
  wire  FA_3_io_cin; // @[RA_Mul.scala 43:21:@3814.4]
  wire  FA_4_io_s; // @[RA_Mul.scala 43:21:@3822.4]
  wire  FA_4_io_cout; // @[RA_Mul.scala 43:21:@3822.4]
  wire  FA_4_io_a; // @[RA_Mul.scala 43:21:@3822.4]
  wire  FA_4_io_b; // @[RA_Mul.scala 43:21:@3822.4]
  wire  FA_4_io_cin; // @[RA_Mul.scala 43:21:@3822.4]
  wire  FA_5_io_s; // @[RA_Mul.scala 43:21:@3830.4]
  wire  FA_5_io_cout; // @[RA_Mul.scala 43:21:@3830.4]
  wire  FA_5_io_a; // @[RA_Mul.scala 43:21:@3830.4]
  wire  FA_5_io_b; // @[RA_Mul.scala 43:21:@3830.4]
  wire  FA_5_io_cin; // @[RA_Mul.scala 43:21:@3830.4]
  wire  FA_6_io_s; // @[RA_Mul.scala 43:21:@3838.4]
  wire  FA_6_io_cout; // @[RA_Mul.scala 43:21:@3838.4]
  wire  FA_6_io_a; // @[RA_Mul.scala 43:21:@3838.4]
  wire  FA_6_io_b; // @[RA_Mul.scala 43:21:@3838.4]
  wire  FA_6_io_cin; // @[RA_Mul.scala 43:21:@3838.4]
  wire  FA_7_io_s; // @[RA_Mul.scala 43:21:@3846.4]
  wire  FA_7_io_cout; // @[RA_Mul.scala 43:21:@3846.4]
  wire  FA_7_io_a; // @[RA_Mul.scala 43:21:@3846.4]
  wire  FA_7_io_b; // @[RA_Mul.scala 43:21:@3846.4]
  wire  FA_7_io_cin; // @[RA_Mul.scala 43:21:@3846.4]
  wire  FA_8_io_s; // @[RA_Mul.scala 43:21:@3854.4]
  wire  FA_8_io_cout; // @[RA_Mul.scala 43:21:@3854.4]
  wire  FA_8_io_a; // @[RA_Mul.scala 43:21:@3854.4]
  wire  FA_8_io_b; // @[RA_Mul.scala 43:21:@3854.4]
  wire  FA_8_io_cin; // @[RA_Mul.scala 43:21:@3854.4]
  wire  FA_9_io_s; // @[RA_Mul.scala 43:21:@3862.4]
  wire  FA_9_io_cout; // @[RA_Mul.scala 43:21:@3862.4]
  wire  FA_9_io_a; // @[RA_Mul.scala 43:21:@3862.4]
  wire  FA_9_io_b; // @[RA_Mul.scala 43:21:@3862.4]
  wire  FA_9_io_cin; // @[RA_Mul.scala 43:21:@3862.4]
  wire  HA_8_io_s; // @[RA_Mul.scala 19:21:@3870.4]
  wire  HA_8_io_cout; // @[RA_Mul.scala 19:21:@3870.4]
  wire  HA_8_io_a; // @[RA_Mul.scala 19:21:@3870.4]
  wire  HA_8_io_b; // @[RA_Mul.scala 19:21:@3870.4]
  wire  FA_10_io_s; // @[RA_Mul.scala 43:21:@3877.4]
  wire  FA_10_io_cout; // @[RA_Mul.scala 43:21:@3877.4]
  wire  FA_10_io_a; // @[RA_Mul.scala 43:21:@3877.4]
  wire  FA_10_io_b; // @[RA_Mul.scala 43:21:@3877.4]
  wire  FA_10_io_cin; // @[RA_Mul.scala 43:21:@3877.4]
  wire  HA_9_io_s; // @[RA_Mul.scala 19:21:@3885.4]
  wire  HA_9_io_cout; // @[RA_Mul.scala 19:21:@3885.4]
  wire  HA_9_io_a; // @[RA_Mul.scala 19:21:@3885.4]
  wire  HA_9_io_b; // @[RA_Mul.scala 19:21:@3885.4]
  wire  FA_11_io_s; // @[RA_Mul.scala 43:21:@3892.4]
  wire  FA_11_io_cout; // @[RA_Mul.scala 43:21:@3892.4]
  wire  FA_11_io_a; // @[RA_Mul.scala 43:21:@3892.4]
  wire  FA_11_io_b; // @[RA_Mul.scala 43:21:@3892.4]
  wire  FA_11_io_cin; // @[RA_Mul.scala 43:21:@3892.4]
  wire  HA_10_io_s; // @[RA_Mul.scala 19:21:@3900.4]
  wire  HA_10_io_cout; // @[RA_Mul.scala 19:21:@3900.4]
  wire  HA_10_io_a; // @[RA_Mul.scala 19:21:@3900.4]
  wire  HA_10_io_b; // @[RA_Mul.scala 19:21:@3900.4]
  wire  FA_12_io_s; // @[RA_Mul.scala 43:21:@3908.4]
  wire  FA_12_io_cout; // @[RA_Mul.scala 43:21:@3908.4]
  wire  FA_12_io_a; // @[RA_Mul.scala 43:21:@3908.4]
  wire  FA_12_io_b; // @[RA_Mul.scala 43:21:@3908.4]
  wire  FA_12_io_cin; // @[RA_Mul.scala 43:21:@3908.4]
  HA HA ( // @[RA_Mul.scala 19:21:@3731.4]
    .io_s(HA_io_s),
    .io_cout(HA_io_cout),
    .io_a(HA_io_a),
    .io_b(HA_io_b)
  );
  FA FA ( // @[RA_Mul.scala 43:21:@3740.4]
    .io_s(FA_io_s),
    .io_cout(FA_io_cout),
    .io_a(FA_io_a),
    .io_b(FA_io_b),
    .io_cin(FA_io_cin)
  );
  HA HA_1 ( // @[RA_Mul.scala 19:21:@3749.4]
    .io_s(HA_1_io_s),
    .io_cout(HA_1_io_cout),
    .io_a(HA_1_io_a),
    .io_b(HA_1_io_b)
  );
  HA HA_2 ( // @[RA_Mul.scala 19:21:@3756.4]
    .io_s(HA_2_io_s),
    .io_cout(HA_2_io_cout),
    .io_a(HA_2_io_a),
    .io_b(HA_2_io_b)
  );
  HA HA_3 ( // @[RA_Mul.scala 19:21:@3763.4]
    .io_s(HA_3_io_s),
    .io_cout(HA_3_io_cout),
    .io_a(HA_3_io_a),
    .io_b(HA_3_io_b)
  );
  HA HA_4 ( // @[RA_Mul.scala 19:21:@3770.4]
    .io_s(HA_4_io_s),
    .io_cout(HA_4_io_cout),
    .io_a(HA_4_io_a),
    .io_b(HA_4_io_b)
  );
  HA HA_5 ( // @[RA_Mul.scala 19:21:@3777.4]
    .io_s(HA_5_io_s),
    .io_cout(HA_5_io_cout),
    .io_a(HA_5_io_a),
    .io_b(HA_5_io_b)
  );
  HA HA_6 ( // @[RA_Mul.scala 19:21:@3784.4]
    .io_s(HA_6_io_s),
    .io_cout(HA_6_io_cout),
    .io_a(HA_6_io_a),
    .io_b(HA_6_io_b)
  );
  HA HA_7 ( // @[RA_Mul.scala 19:21:@3791.4]
    .io_s(HA_7_io_s),
    .io_cout(HA_7_io_cout),
    .io_a(HA_7_io_a),
    .io_b(HA_7_io_b)
  );
  FA FA_1 ( // @[RA_Mul.scala 43:21:@3798.4]
    .io_s(FA_1_io_s),
    .io_cout(FA_1_io_cout),
    .io_a(FA_1_io_a),
    .io_b(FA_1_io_b),
    .io_cin(FA_1_io_cin)
  );
  FA FA_2 ( // @[RA_Mul.scala 43:21:@3806.4]
    .io_s(FA_2_io_s),
    .io_cout(FA_2_io_cout),
    .io_a(FA_2_io_a),
    .io_b(FA_2_io_b),
    .io_cin(FA_2_io_cin)
  );
  FA FA_3 ( // @[RA_Mul.scala 43:21:@3814.4]
    .io_s(FA_3_io_s),
    .io_cout(FA_3_io_cout),
    .io_a(FA_3_io_a),
    .io_b(FA_3_io_b),
    .io_cin(FA_3_io_cin)
  );
  FA FA_4 ( // @[RA_Mul.scala 43:21:@3822.4]
    .io_s(FA_4_io_s),
    .io_cout(FA_4_io_cout),
    .io_a(FA_4_io_a),
    .io_b(FA_4_io_b),
    .io_cin(FA_4_io_cin)
  );
  FA FA_5 ( // @[RA_Mul.scala 43:21:@3830.4]
    .io_s(FA_5_io_s),
    .io_cout(FA_5_io_cout),
    .io_a(FA_5_io_a),
    .io_b(FA_5_io_b),
    .io_cin(FA_5_io_cin)
  );
  FA FA_6 ( // @[RA_Mul.scala 43:21:@3838.4]
    .io_s(FA_6_io_s),
    .io_cout(FA_6_io_cout),
    .io_a(FA_6_io_a),
    .io_b(FA_6_io_b),
    .io_cin(FA_6_io_cin)
  );
  FA FA_7 ( // @[RA_Mul.scala 43:21:@3846.4]
    .io_s(FA_7_io_s),
    .io_cout(FA_7_io_cout),
    .io_a(FA_7_io_a),
    .io_b(FA_7_io_b),
    .io_cin(FA_7_io_cin)
  );
  FA FA_8 ( // @[RA_Mul.scala 43:21:@3854.4]
    .io_s(FA_8_io_s),
    .io_cout(FA_8_io_cout),
    .io_a(FA_8_io_a),
    .io_b(FA_8_io_b),
    .io_cin(FA_8_io_cin)
  );
  FA FA_9 ( // @[RA_Mul.scala 43:21:@3862.4]
    .io_s(FA_9_io_s),
    .io_cout(FA_9_io_cout),
    .io_a(FA_9_io_a),
    .io_b(FA_9_io_b),
    .io_cin(FA_9_io_cin)
  );
  HA HA_8 ( // @[RA_Mul.scala 19:21:@3870.4]
    .io_s(HA_8_io_s),
    .io_cout(HA_8_io_cout),
    .io_a(HA_8_io_a),
    .io_b(HA_8_io_b)
  );
  FA FA_10 ( // @[RA_Mul.scala 43:21:@3877.4]
    .io_s(FA_10_io_s),
    .io_cout(FA_10_io_cout),
    .io_a(FA_10_io_a),
    .io_b(FA_10_io_b),
    .io_cin(FA_10_io_cin)
  );
  HA HA_9 ( // @[RA_Mul.scala 19:21:@3885.4]
    .io_s(HA_9_io_s),
    .io_cout(HA_9_io_cout),
    .io_a(HA_9_io_a),
    .io_b(HA_9_io_b)
  );
  FA FA_11 ( // @[RA_Mul.scala 43:21:@3892.4]
    .io_s(FA_11_io_s),
    .io_cout(FA_11_io_cout),
    .io_a(FA_11_io_a),
    .io_b(FA_11_io_b),
    .io_cin(FA_11_io_cin)
  );
  HA HA_10 ( // @[RA_Mul.scala 19:21:@3900.4]
    .io_s(HA_10_io_s),
    .io_cout(HA_10_io_cout),
    .io_a(HA_10_io_a),
    .io_b(HA_10_io_b)
  );
  FA FA_12 ( // @[RA_Mul.scala 43:21:@3908.4]
    .io_s(FA_12_io_s),
    .io_cout(FA_12_io_cout),
    .io_a(FA_12_io_a),
    .io_b(FA_12_io_b),
    .io_cin(FA_12_io_cin)
  );
  assign io_matrix_o_0_0 = io_matrix_i_0_0; // @[RA_Mul.scala 555:23:@3725.4]
  assign io_matrix_o_0_1 = io_matrix_i_0_1; // @[RA_Mul.scala 555:23:@3727.4]
  assign io_matrix_o_0_2 = io_matrix_i_0_2; // @[RA_Mul.scala 555:23:@3729.4]
  assign io_matrix_o_0_3 = HA_io_s; // @[RA_Mul.scala 22:7:@3736.4]
  assign io_matrix_o_0_4 = io_matrix_i_0_4; // @[RA_Mul.scala 562:21:@3739.4]
  assign io_matrix_o_0_5 = FA_io_s; // @[RA_Mul.scala 47:7:@3746.4]
  assign io_matrix_o_0_6 = HA_1_io_s; // @[RA_Mul.scala 22:7:@3754.4]
  assign io_matrix_o_0_7 = HA_2_io_s; // @[RA_Mul.scala 22:7:@3761.4]
  assign io_matrix_o_0_8 = HA_3_io_s; // @[RA_Mul.scala 22:7:@3768.4]
  assign io_matrix_o_0_9 = HA_4_io_s; // @[RA_Mul.scala 22:7:@3775.4]
  assign io_matrix_o_0_10 = HA_5_io_s; // @[RA_Mul.scala 22:7:@3782.4]
  assign io_matrix_o_0_11 = HA_6_io_s; // @[RA_Mul.scala 22:7:@3789.4]
  assign io_matrix_o_0_12 = HA_7_io_s; // @[RA_Mul.scala 22:7:@3796.4]
  assign io_matrix_o_0_13 = FA_1_io_s; // @[RA_Mul.scala 47:7:@3804.4]
  assign io_matrix_o_0_14 = FA_2_io_s; // @[RA_Mul.scala 47:7:@3812.4]
  assign io_matrix_o_0_15 = FA_3_io_s; // @[RA_Mul.scala 47:7:@3820.4]
  assign io_matrix_o_0_16 = FA_4_io_s; // @[RA_Mul.scala 47:7:@3828.4]
  assign io_matrix_o_0_17 = FA_5_io_s; // @[RA_Mul.scala 47:7:@3836.4]
  assign io_matrix_o_0_18 = FA_6_io_s; // @[RA_Mul.scala 47:7:@3844.4]
  assign io_matrix_o_0_19 = FA_7_io_s; // @[RA_Mul.scala 47:7:@3852.4]
  assign io_matrix_o_0_20 = FA_8_io_s; // @[RA_Mul.scala 47:7:@3860.4]
  assign io_matrix_o_0_21 = FA_9_io_s; // @[RA_Mul.scala 47:7:@3868.4]
  assign io_matrix_o_0_22 = HA_8_io_s; // @[RA_Mul.scala 22:7:@3875.4]
  assign io_matrix_o_0_23 = FA_10_io_s; // @[RA_Mul.scala 47:7:@3883.4]
  assign io_matrix_o_0_24 = HA_9_io_s; // @[RA_Mul.scala 22:7:@3890.4]
  assign io_matrix_o_0_25 = FA_11_io_s; // @[RA_Mul.scala 47:7:@3898.4]
  assign io_matrix_o_0_26 = HA_10_io_s; // @[RA_Mul.scala 22:7:@3905.4]
  assign io_matrix_o_0_27 = io_matrix_i_0_27; // @[RA_Mul.scala 582:22:@3907.4]
  assign io_matrix_o_0_28 = FA_12_io_s; // @[RA_Mul.scala 47:7:@3914.4]
  assign io_matrix_o_0_29 = io_matrix_i_0_29; // @[RA_Mul.scala 587:22:@3917.4]
  assign io_matrix_o_0_30 = io_matrix_i_0_30; // @[RA_Mul.scala 589:22:@3918.4]
  assign io_matrix_o_0_31 = io_matrix_i_0_31; // @[RA_Mul.scala 592:22:@3920.4]
  assign io_matrix_o_1_4 = HA_io_cout; // @[RA_Mul.scala 23:10:@3737.4]
  assign io_matrix_o_1_6 = FA_io_cout; // @[RA_Mul.scala 48:10:@3747.4]
  assign io_matrix_o_1_7 = HA_1_io_cout; // @[RA_Mul.scala 23:10:@3755.4]
  assign io_matrix_o_1_8 = HA_2_io_cout; // @[RA_Mul.scala 23:10:@3762.4]
  assign io_matrix_o_1_9 = HA_3_io_cout; // @[RA_Mul.scala 23:10:@3769.4]
  assign io_matrix_o_1_10 = HA_4_io_cout; // @[RA_Mul.scala 23:10:@3776.4]
  assign io_matrix_o_1_11 = HA_5_io_cout; // @[RA_Mul.scala 23:10:@3783.4]
  assign io_matrix_o_1_12 = HA_6_io_cout; // @[RA_Mul.scala 23:10:@3790.4]
  assign io_matrix_o_1_13 = HA_7_io_cout; // @[RA_Mul.scala 23:10:@3797.4]
  assign io_matrix_o_1_14 = FA_1_io_cout; // @[RA_Mul.scala 48:10:@3805.4]
  assign io_matrix_o_1_15 = FA_2_io_cout; // @[RA_Mul.scala 48:10:@3813.4]
  assign io_matrix_o_1_16 = FA_3_io_cout; // @[RA_Mul.scala 48:10:@3821.4]
  assign io_matrix_o_1_17 = FA_4_io_cout; // @[RA_Mul.scala 48:10:@3829.4]
  assign io_matrix_o_1_18 = FA_5_io_cout; // @[RA_Mul.scala 48:10:@3837.4]
  assign io_matrix_o_1_19 = FA_6_io_cout; // @[RA_Mul.scala 48:10:@3845.4]
  assign io_matrix_o_1_20 = FA_7_io_cout; // @[RA_Mul.scala 48:10:@3853.4]
  assign io_matrix_o_1_21 = FA_8_io_cout; // @[RA_Mul.scala 48:10:@3861.4]
  assign io_matrix_o_1_22 = FA_9_io_cout; // @[RA_Mul.scala 48:10:@3869.4]
  assign io_matrix_o_1_23 = HA_8_io_cout; // @[RA_Mul.scala 23:10:@3876.4]
  assign io_matrix_o_1_24 = FA_10_io_cout; // @[RA_Mul.scala 48:10:@3884.4]
  assign io_matrix_o_1_25 = HA_9_io_cout; // @[RA_Mul.scala 23:10:@3891.4]
  assign io_matrix_o_1_26 = FA_11_io_cout; // @[RA_Mul.scala 48:10:@3899.4]
  assign io_matrix_o_1_27 = HA_10_io_cout; // @[RA_Mul.scala 23:10:@3906.4]
  assign io_matrix_o_1_29 = FA_12_io_cout; // @[RA_Mul.scala 48:10:@3915.4]
  assign io_matrix_o_1_31 = io_matrix_i_1_31; // @[RA_Mul.scala 593:22:@3921.4]
  assign HA_io_a = io_matrix_i_0_3; // @[RA_Mul.scala 20:14:@3734.4]
  assign HA_io_b = io_matrix_i_1_3; // @[RA_Mul.scala 21:14:@3735.4]
  assign FA_io_a = io_matrix_i_0_5; // @[RA_Mul.scala 44:14:@3743.4]
  assign FA_io_b = io_matrix_i_1_5; // @[RA_Mul.scala 45:14:@3744.4]
  assign FA_io_cin = io_matrix_i_2_5; // @[RA_Mul.scala 46:16:@3745.4]
  assign HA_1_io_a = io_matrix_i_0_6; // @[RA_Mul.scala 20:14:@3752.4]
  assign HA_1_io_b = io_matrix_i_1_6; // @[RA_Mul.scala 21:14:@3753.4]
  assign HA_2_io_a = io_matrix_i_0_7; // @[RA_Mul.scala 20:14:@3759.4]
  assign HA_2_io_b = io_matrix_i_1_7; // @[RA_Mul.scala 21:14:@3760.4]
  assign HA_3_io_a = io_matrix_i_0_8; // @[RA_Mul.scala 20:14:@3766.4]
  assign HA_3_io_b = io_matrix_i_1_8; // @[RA_Mul.scala 21:14:@3767.4]
  assign HA_4_io_a = io_matrix_i_0_9; // @[RA_Mul.scala 20:14:@3773.4]
  assign HA_4_io_b = io_matrix_i_1_9; // @[RA_Mul.scala 21:14:@3774.4]
  assign HA_5_io_a = io_matrix_i_0_10; // @[RA_Mul.scala 20:14:@3780.4]
  assign HA_5_io_b = io_matrix_i_1_10; // @[RA_Mul.scala 21:14:@3781.4]
  assign HA_6_io_a = io_matrix_i_0_11; // @[RA_Mul.scala 20:14:@3787.4]
  assign HA_6_io_b = io_matrix_i_1_11; // @[RA_Mul.scala 21:14:@3788.4]
  assign HA_7_io_a = io_matrix_i_0_12; // @[RA_Mul.scala 20:14:@3794.4]
  assign HA_7_io_b = io_matrix_i_1_12; // @[RA_Mul.scala 21:14:@3795.4]
  assign FA_1_io_a = io_matrix_i_0_13; // @[RA_Mul.scala 44:14:@3801.4]
  assign FA_1_io_b = io_matrix_i_1_13; // @[RA_Mul.scala 45:14:@3802.4]
  assign FA_1_io_cin = io_matrix_i_2_13; // @[RA_Mul.scala 46:16:@3803.4]
  assign FA_2_io_a = io_matrix_i_0_14; // @[RA_Mul.scala 44:14:@3809.4]
  assign FA_2_io_b = io_matrix_i_1_14; // @[RA_Mul.scala 45:14:@3810.4]
  assign FA_2_io_cin = io_matrix_i_2_14; // @[RA_Mul.scala 46:16:@3811.4]
  assign FA_3_io_a = io_matrix_i_0_15; // @[RA_Mul.scala 44:14:@3817.4]
  assign FA_3_io_b = io_matrix_i_1_15; // @[RA_Mul.scala 45:14:@3818.4]
  assign FA_3_io_cin = io_matrix_i_2_15; // @[RA_Mul.scala 46:16:@3819.4]
  assign FA_4_io_a = io_matrix_i_0_16; // @[RA_Mul.scala 44:14:@3825.4]
  assign FA_4_io_b = io_matrix_i_1_16; // @[RA_Mul.scala 45:14:@3826.4]
  assign FA_4_io_cin = io_matrix_i_2_16; // @[RA_Mul.scala 46:16:@3827.4]
  assign FA_5_io_a = io_matrix_i_0_17; // @[RA_Mul.scala 44:14:@3833.4]
  assign FA_5_io_b = io_matrix_i_1_17; // @[RA_Mul.scala 45:14:@3834.4]
  assign FA_5_io_cin = io_matrix_i_2_17; // @[RA_Mul.scala 46:16:@3835.4]
  assign FA_6_io_a = io_matrix_i_0_18; // @[RA_Mul.scala 44:14:@3841.4]
  assign FA_6_io_b = io_matrix_i_1_18; // @[RA_Mul.scala 45:14:@3842.4]
  assign FA_6_io_cin = io_matrix_i_2_18; // @[RA_Mul.scala 46:16:@3843.4]
  assign FA_7_io_a = io_matrix_i_0_19; // @[RA_Mul.scala 44:14:@3849.4]
  assign FA_7_io_b = io_matrix_i_1_19; // @[RA_Mul.scala 45:14:@3850.4]
  assign FA_7_io_cin = io_matrix_i_2_19; // @[RA_Mul.scala 46:16:@3851.4]
  assign FA_8_io_a = io_matrix_i_0_20; // @[RA_Mul.scala 44:14:@3857.4]
  assign FA_8_io_b = io_matrix_i_1_20; // @[RA_Mul.scala 45:14:@3858.4]
  assign FA_8_io_cin = io_matrix_i_2_20; // @[RA_Mul.scala 46:16:@3859.4]
  assign FA_9_io_a = io_matrix_i_0_21; // @[RA_Mul.scala 44:14:@3865.4]
  assign FA_9_io_b = io_matrix_i_1_21; // @[RA_Mul.scala 45:14:@3866.4]
  assign FA_9_io_cin = io_matrix_i_2_21; // @[RA_Mul.scala 46:16:@3867.4]
  assign HA_8_io_a = io_matrix_i_0_22; // @[RA_Mul.scala 20:14:@3873.4]
  assign HA_8_io_b = io_matrix_i_1_22; // @[RA_Mul.scala 21:14:@3874.4]
  assign FA_10_io_a = io_matrix_i_0_23; // @[RA_Mul.scala 44:14:@3880.4]
  assign FA_10_io_b = io_matrix_i_1_23; // @[RA_Mul.scala 45:14:@3881.4]
  assign FA_10_io_cin = io_matrix_i_2_23; // @[RA_Mul.scala 46:16:@3882.4]
  assign HA_9_io_a = io_matrix_i_0_24; // @[RA_Mul.scala 20:14:@3888.4]
  assign HA_9_io_b = io_matrix_i_1_24; // @[RA_Mul.scala 21:14:@3889.4]
  assign FA_11_io_a = io_matrix_i_0_25; // @[RA_Mul.scala 44:14:@3895.4]
  assign FA_11_io_b = io_matrix_i_1_25; // @[RA_Mul.scala 45:14:@3896.4]
  assign FA_11_io_cin = io_matrix_i_2_25; // @[RA_Mul.scala 46:16:@3897.4]
  assign HA_10_io_a = io_matrix_i_0_26; // @[RA_Mul.scala 20:14:@3903.4]
  assign HA_10_io_b = io_matrix_i_1_26; // @[RA_Mul.scala 21:14:@3904.4]
  assign FA_12_io_a = io_matrix_i_0_28; // @[RA_Mul.scala 44:14:@3911.4]
  assign FA_12_io_b = io_matrix_i_1_28; // @[RA_Mul.scala 45:14:@3912.4]
  assign FA_12_io_cin = io_matrix_i_2_28; // @[RA_Mul.scala 46:16:@3913.4]
endmodule
module PPLRegs2( // @[:@3923.2]
  input   clock, // @[:@3924.4]
  input   reset, // @[:@3925.4]
  output  io_matrix_o_0_0, // @[:@3926.4]
  output  io_matrix_o_0_1, // @[:@3926.4]
  output  io_matrix_o_0_2, // @[:@3926.4]
  output  io_matrix_o_0_3, // @[:@3926.4]
  output  io_matrix_o_0_4, // @[:@3926.4]
  output  io_matrix_o_0_5, // @[:@3926.4]
  output  io_matrix_o_0_6, // @[:@3926.4]
  output  io_matrix_o_0_7, // @[:@3926.4]
  output  io_matrix_o_0_8, // @[:@3926.4]
  output  io_matrix_o_0_9, // @[:@3926.4]
  output  io_matrix_o_0_10, // @[:@3926.4]
  output  io_matrix_o_0_11, // @[:@3926.4]
  output  io_matrix_o_0_12, // @[:@3926.4]
  output  io_matrix_o_0_13, // @[:@3926.4]
  output  io_matrix_o_0_14, // @[:@3926.4]
  output  io_matrix_o_0_15, // @[:@3926.4]
  output  io_matrix_o_0_16, // @[:@3926.4]
  output  io_matrix_o_0_17, // @[:@3926.4]
  output  io_matrix_o_0_18, // @[:@3926.4]
  output  io_matrix_o_0_19, // @[:@3926.4]
  output  io_matrix_o_0_20, // @[:@3926.4]
  output  io_matrix_o_0_21, // @[:@3926.4]
  output  io_matrix_o_0_22, // @[:@3926.4]
  output  io_matrix_o_0_23, // @[:@3926.4]
  output  io_matrix_o_0_24, // @[:@3926.4]
  output  io_matrix_o_0_25, // @[:@3926.4]
  output  io_matrix_o_0_26, // @[:@3926.4]
  output  io_matrix_o_0_27, // @[:@3926.4]
  output  io_matrix_o_0_28, // @[:@3926.4]
  output  io_matrix_o_0_29, // @[:@3926.4]
  output  io_matrix_o_0_30, // @[:@3926.4]
  output  io_matrix_o_0_31, // @[:@3926.4]
  output  io_matrix_o_1_0, // @[:@3926.4]
  output  io_matrix_o_1_1, // @[:@3926.4]
  output  io_matrix_o_1_2, // @[:@3926.4]
  output  io_matrix_o_1_3, // @[:@3926.4]
  output  io_matrix_o_1_4, // @[:@3926.4]
  output  io_matrix_o_1_5, // @[:@3926.4]
  output  io_matrix_o_1_6, // @[:@3926.4]
  output  io_matrix_o_1_7, // @[:@3926.4]
  output  io_matrix_o_1_8, // @[:@3926.4]
  output  io_matrix_o_1_9, // @[:@3926.4]
  output  io_matrix_o_1_10, // @[:@3926.4]
  output  io_matrix_o_1_11, // @[:@3926.4]
  output  io_matrix_o_1_12, // @[:@3926.4]
  output  io_matrix_o_1_13, // @[:@3926.4]
  output  io_matrix_o_1_14, // @[:@3926.4]
  output  io_matrix_o_1_15, // @[:@3926.4]
  output  io_matrix_o_1_16, // @[:@3926.4]
  output  io_matrix_o_1_17, // @[:@3926.4]
  output  io_matrix_o_1_18, // @[:@3926.4]
  output  io_matrix_o_1_19, // @[:@3926.4]
  output  io_matrix_o_1_20, // @[:@3926.4]
  output  io_matrix_o_1_21, // @[:@3926.4]
  output  io_matrix_o_1_22, // @[:@3926.4]
  output  io_matrix_o_1_23, // @[:@3926.4]
  output  io_matrix_o_1_24, // @[:@3926.4]
  output  io_matrix_o_1_25, // @[:@3926.4]
  output  io_matrix_o_1_26, // @[:@3926.4]
  output  io_matrix_o_1_27, // @[:@3926.4]
  output  io_matrix_o_1_28, // @[:@3926.4]
  output  io_matrix_o_1_29, // @[:@3926.4]
  output  io_matrix_o_1_30, // @[:@3926.4]
  output  io_matrix_o_1_31, // @[:@3926.4]
  input   io_matrix_i_0_0, // @[:@3926.4]
  input   io_matrix_i_0_1, // @[:@3926.4]
  input   io_matrix_i_0_2, // @[:@3926.4]
  input   io_matrix_i_0_3, // @[:@3926.4]
  input   io_matrix_i_0_4, // @[:@3926.4]
  input   io_matrix_i_0_5, // @[:@3926.4]
  input   io_matrix_i_0_6, // @[:@3926.4]
  input   io_matrix_i_0_7, // @[:@3926.4]
  input   io_matrix_i_0_8, // @[:@3926.4]
  input   io_matrix_i_0_9, // @[:@3926.4]
  input   io_matrix_i_0_10, // @[:@3926.4]
  input   io_matrix_i_0_11, // @[:@3926.4]
  input   io_matrix_i_0_12, // @[:@3926.4]
  input   io_matrix_i_0_13, // @[:@3926.4]
  input   io_matrix_i_0_14, // @[:@3926.4]
  input   io_matrix_i_0_15, // @[:@3926.4]
  input   io_matrix_i_0_16, // @[:@3926.4]
  input   io_matrix_i_0_17, // @[:@3926.4]
  input   io_matrix_i_0_18, // @[:@3926.4]
  input   io_matrix_i_0_19, // @[:@3926.4]
  input   io_matrix_i_0_20, // @[:@3926.4]
  input   io_matrix_i_0_21, // @[:@3926.4]
  input   io_matrix_i_0_22, // @[:@3926.4]
  input   io_matrix_i_0_23, // @[:@3926.4]
  input   io_matrix_i_0_24, // @[:@3926.4]
  input   io_matrix_i_0_25, // @[:@3926.4]
  input   io_matrix_i_0_26, // @[:@3926.4]
  input   io_matrix_i_0_27, // @[:@3926.4]
  input   io_matrix_i_0_28, // @[:@3926.4]
  input   io_matrix_i_0_29, // @[:@3926.4]
  input   io_matrix_i_0_30, // @[:@3926.4]
  input   io_matrix_i_0_31, // @[:@3926.4]
  input   io_matrix_i_1_4, // @[:@3926.4]
  input   io_matrix_i_1_6, // @[:@3926.4]
  input   io_matrix_i_1_7, // @[:@3926.4]
  input   io_matrix_i_1_8, // @[:@3926.4]
  input   io_matrix_i_1_9, // @[:@3926.4]
  input   io_matrix_i_1_10, // @[:@3926.4]
  input   io_matrix_i_1_11, // @[:@3926.4]
  input   io_matrix_i_1_12, // @[:@3926.4]
  input   io_matrix_i_1_13, // @[:@3926.4]
  input   io_matrix_i_1_14, // @[:@3926.4]
  input   io_matrix_i_1_15, // @[:@3926.4]
  input   io_matrix_i_1_16, // @[:@3926.4]
  input   io_matrix_i_1_17, // @[:@3926.4]
  input   io_matrix_i_1_18, // @[:@3926.4]
  input   io_matrix_i_1_19, // @[:@3926.4]
  input   io_matrix_i_1_20, // @[:@3926.4]
  input   io_matrix_i_1_21, // @[:@3926.4]
  input   io_matrix_i_1_22, // @[:@3926.4]
  input   io_matrix_i_1_23, // @[:@3926.4]
  input   io_matrix_i_1_24, // @[:@3926.4]
  input   io_matrix_i_1_25, // @[:@3926.4]
  input   io_matrix_i_1_26, // @[:@3926.4]
  input   io_matrix_i_1_27, // @[:@3926.4]
  input   io_matrix_i_1_29, // @[:@3926.4]
  input   io_matrix_i_1_31 // @[:@3926.4]
);
  wire [1:0] _T_1668; // @[RA_Mul.scala 702:21:@3929.4]
  wire [1:0] _T_1669; // @[RA_Mul.scala 702:21:@3930.4]
  wire [3:0] _T_1670; // @[RA_Mul.scala 702:21:@3931.4]
  wire [1:0] _T_1671; // @[RA_Mul.scala 702:21:@3932.4]
  wire [1:0] _T_1672; // @[RA_Mul.scala 702:21:@3933.4]
  wire [3:0] _T_1673; // @[RA_Mul.scala 702:21:@3934.4]
  wire [7:0] _T_1674; // @[RA_Mul.scala 702:21:@3935.4]
  wire [1:0] _T_1675; // @[RA_Mul.scala 702:21:@3936.4]
  wire [1:0] _T_1676; // @[RA_Mul.scala 702:21:@3937.4]
  wire [3:0] _T_1677; // @[RA_Mul.scala 702:21:@3938.4]
  wire [1:0] _T_1678; // @[RA_Mul.scala 702:21:@3939.4]
  wire [1:0] _T_1679; // @[RA_Mul.scala 702:21:@3940.4]
  wire [3:0] _T_1680; // @[RA_Mul.scala 702:21:@3941.4]
  wire [7:0] _T_1681; // @[RA_Mul.scala 702:21:@3942.4]
  wire [15:0] _T_1682; // @[RA_Mul.scala 702:21:@3943.4]
  wire [1:0] _T_1683; // @[RA_Mul.scala 702:21:@3944.4]
  wire [1:0] _T_1684; // @[RA_Mul.scala 702:21:@3945.4]
  wire [3:0] _T_1685; // @[RA_Mul.scala 702:21:@3946.4]
  wire [1:0] _T_1686; // @[RA_Mul.scala 702:21:@3947.4]
  wire [1:0] _T_1687; // @[RA_Mul.scala 702:21:@3948.4]
  wire [3:0] _T_1688; // @[RA_Mul.scala 702:21:@3949.4]
  wire [7:0] _T_1689; // @[RA_Mul.scala 702:21:@3950.4]
  wire [1:0] _T_1690; // @[RA_Mul.scala 702:21:@3951.4]
  wire [1:0] _T_1691; // @[RA_Mul.scala 702:21:@3952.4]
  wire [3:0] _T_1692; // @[RA_Mul.scala 702:21:@3953.4]
  wire [1:0] _T_1693; // @[RA_Mul.scala 702:21:@3954.4]
  wire [1:0] _T_1694; // @[RA_Mul.scala 702:21:@3955.4]
  wire [3:0] _T_1695; // @[RA_Mul.scala 702:21:@3956.4]
  wire [7:0] _T_1696; // @[RA_Mul.scala 702:21:@3957.4]
  wire [15:0] _T_1697; // @[RA_Mul.scala 702:21:@3958.4]
  wire [31:0] _T_1698; // @[RA_Mul.scala 702:21:@3959.4]
  reg [31:0] tmp_0; // @[RA_Mul.scala 702:18:@3960.4]
  reg [31:0] _RAND_0;
  wire [1:0] _T_1705; // @[RA_Mul.scala 702:21:@3966.4]
  wire [1:0] _T_1706; // @[RA_Mul.scala 702:21:@3967.4]
  wire [3:0] _T_1707; // @[RA_Mul.scala 702:21:@3968.4]
  wire [7:0] _T_1708; // @[RA_Mul.scala 702:21:@3969.4]
  wire [1:0] _T_1709; // @[RA_Mul.scala 702:21:@3970.4]
  wire [1:0] _T_1710; // @[RA_Mul.scala 702:21:@3971.4]
  wire [3:0] _T_1711; // @[RA_Mul.scala 702:21:@3972.4]
  wire [1:0] _T_1712; // @[RA_Mul.scala 702:21:@3973.4]
  wire [1:0] _T_1713; // @[RA_Mul.scala 702:21:@3974.4]
  wire [3:0] _T_1714; // @[RA_Mul.scala 702:21:@3975.4]
  wire [7:0] _T_1715; // @[RA_Mul.scala 702:21:@3976.4]
  wire [15:0] _T_1716; // @[RA_Mul.scala 702:21:@3977.4]
  wire [1:0] _T_1717; // @[RA_Mul.scala 702:21:@3978.4]
  wire [1:0] _T_1718; // @[RA_Mul.scala 702:21:@3979.4]
  wire [3:0] _T_1719; // @[RA_Mul.scala 702:21:@3980.4]
  wire [1:0] _T_1720; // @[RA_Mul.scala 702:21:@3981.4]
  wire [1:0] _T_1721; // @[RA_Mul.scala 702:21:@3982.4]
  wire [3:0] _T_1722; // @[RA_Mul.scala 702:21:@3983.4]
  wire [7:0] _T_1723; // @[RA_Mul.scala 702:21:@3984.4]
  wire [1:0] _T_1724; // @[RA_Mul.scala 702:21:@3985.4]
  wire [1:0] _T_1725; // @[RA_Mul.scala 702:21:@3986.4]
  wire [3:0] _T_1726; // @[RA_Mul.scala 702:21:@3987.4]
  wire [1:0] _T_1727; // @[RA_Mul.scala 702:21:@3988.4]
  wire [1:0] _T_1728; // @[RA_Mul.scala 702:21:@3989.4]
  wire [3:0] _T_1729; // @[RA_Mul.scala 702:21:@3990.4]
  wire [7:0] _T_1730; // @[RA_Mul.scala 702:21:@3991.4]
  wire [15:0] _T_1731; // @[RA_Mul.scala 702:21:@3992.4]
  wire [31:0] _T_1732; // @[RA_Mul.scala 702:21:@3993.4]
  reg [31:0] tmp_1; // @[RA_Mul.scala 702:18:@3994.4]
  reg [31:0] _RAND_1;
  assign _T_1668 = {io_matrix_i_0_1,io_matrix_i_0_0}; // @[RA_Mul.scala 702:21:@3929.4]
  assign _T_1669 = {io_matrix_i_0_3,io_matrix_i_0_2}; // @[RA_Mul.scala 702:21:@3930.4]
  assign _T_1670 = {_T_1669,_T_1668}; // @[RA_Mul.scala 702:21:@3931.4]
  assign _T_1671 = {io_matrix_i_0_5,io_matrix_i_0_4}; // @[RA_Mul.scala 702:21:@3932.4]
  assign _T_1672 = {io_matrix_i_0_7,io_matrix_i_0_6}; // @[RA_Mul.scala 702:21:@3933.4]
  assign _T_1673 = {_T_1672,_T_1671}; // @[RA_Mul.scala 702:21:@3934.4]
  assign _T_1674 = {_T_1673,_T_1670}; // @[RA_Mul.scala 702:21:@3935.4]
  assign _T_1675 = {io_matrix_i_0_9,io_matrix_i_0_8}; // @[RA_Mul.scala 702:21:@3936.4]
  assign _T_1676 = {io_matrix_i_0_11,io_matrix_i_0_10}; // @[RA_Mul.scala 702:21:@3937.4]
  assign _T_1677 = {_T_1676,_T_1675}; // @[RA_Mul.scala 702:21:@3938.4]
  assign _T_1678 = {io_matrix_i_0_13,io_matrix_i_0_12}; // @[RA_Mul.scala 702:21:@3939.4]
  assign _T_1679 = {io_matrix_i_0_15,io_matrix_i_0_14}; // @[RA_Mul.scala 702:21:@3940.4]
  assign _T_1680 = {_T_1679,_T_1678}; // @[RA_Mul.scala 702:21:@3941.4]
  assign _T_1681 = {_T_1680,_T_1677}; // @[RA_Mul.scala 702:21:@3942.4]
  assign _T_1682 = {_T_1681,_T_1674}; // @[RA_Mul.scala 702:21:@3943.4]
  assign _T_1683 = {io_matrix_i_0_17,io_matrix_i_0_16}; // @[RA_Mul.scala 702:21:@3944.4]
  assign _T_1684 = {io_matrix_i_0_19,io_matrix_i_0_18}; // @[RA_Mul.scala 702:21:@3945.4]
  assign _T_1685 = {_T_1684,_T_1683}; // @[RA_Mul.scala 702:21:@3946.4]
  assign _T_1686 = {io_matrix_i_0_21,io_matrix_i_0_20}; // @[RA_Mul.scala 702:21:@3947.4]
  assign _T_1687 = {io_matrix_i_0_23,io_matrix_i_0_22}; // @[RA_Mul.scala 702:21:@3948.4]
  assign _T_1688 = {_T_1687,_T_1686}; // @[RA_Mul.scala 702:21:@3949.4]
  assign _T_1689 = {_T_1688,_T_1685}; // @[RA_Mul.scala 702:21:@3950.4]
  assign _T_1690 = {io_matrix_i_0_25,io_matrix_i_0_24}; // @[RA_Mul.scala 702:21:@3951.4]
  assign _T_1691 = {io_matrix_i_0_27,io_matrix_i_0_26}; // @[RA_Mul.scala 702:21:@3952.4]
  assign _T_1692 = {_T_1691,_T_1690}; // @[RA_Mul.scala 702:21:@3953.4]
  assign _T_1693 = {io_matrix_i_0_29,io_matrix_i_0_28}; // @[RA_Mul.scala 702:21:@3954.4]
  assign _T_1694 = {io_matrix_i_0_31,io_matrix_i_0_30}; // @[RA_Mul.scala 702:21:@3955.4]
  assign _T_1695 = {_T_1694,_T_1693}; // @[RA_Mul.scala 702:21:@3956.4]
  assign _T_1696 = {_T_1695,_T_1692}; // @[RA_Mul.scala 702:21:@3957.4]
  assign _T_1697 = {_T_1696,_T_1689}; // @[RA_Mul.scala 702:21:@3958.4]
  assign _T_1698 = {_T_1697,_T_1682}; // @[RA_Mul.scala 702:21:@3959.4]
  assign _T_1705 = {1'h0,io_matrix_i_1_4}; // @[RA_Mul.scala 702:21:@3966.4]
  assign _T_1706 = {io_matrix_i_1_7,io_matrix_i_1_6}; // @[RA_Mul.scala 702:21:@3967.4]
  assign _T_1707 = {_T_1706,_T_1705}; // @[RA_Mul.scala 702:21:@3968.4]
  assign _T_1708 = {_T_1707,4'h0}; // @[RA_Mul.scala 702:21:@3969.4]
  assign _T_1709 = {io_matrix_i_1_9,io_matrix_i_1_8}; // @[RA_Mul.scala 702:21:@3970.4]
  assign _T_1710 = {io_matrix_i_1_11,io_matrix_i_1_10}; // @[RA_Mul.scala 702:21:@3971.4]
  assign _T_1711 = {_T_1710,_T_1709}; // @[RA_Mul.scala 702:21:@3972.4]
  assign _T_1712 = {io_matrix_i_1_13,io_matrix_i_1_12}; // @[RA_Mul.scala 702:21:@3973.4]
  assign _T_1713 = {io_matrix_i_1_15,io_matrix_i_1_14}; // @[RA_Mul.scala 702:21:@3974.4]
  assign _T_1714 = {_T_1713,_T_1712}; // @[RA_Mul.scala 702:21:@3975.4]
  assign _T_1715 = {_T_1714,_T_1711}; // @[RA_Mul.scala 702:21:@3976.4]
  assign _T_1716 = {_T_1715,_T_1708}; // @[RA_Mul.scala 702:21:@3977.4]
  assign _T_1717 = {io_matrix_i_1_17,io_matrix_i_1_16}; // @[RA_Mul.scala 702:21:@3978.4]
  assign _T_1718 = {io_matrix_i_1_19,io_matrix_i_1_18}; // @[RA_Mul.scala 702:21:@3979.4]
  assign _T_1719 = {_T_1718,_T_1717}; // @[RA_Mul.scala 702:21:@3980.4]
  assign _T_1720 = {io_matrix_i_1_21,io_matrix_i_1_20}; // @[RA_Mul.scala 702:21:@3981.4]
  assign _T_1721 = {io_matrix_i_1_23,io_matrix_i_1_22}; // @[RA_Mul.scala 702:21:@3982.4]
  assign _T_1722 = {_T_1721,_T_1720}; // @[RA_Mul.scala 702:21:@3983.4]
  assign _T_1723 = {_T_1722,_T_1719}; // @[RA_Mul.scala 702:21:@3984.4]
  assign _T_1724 = {io_matrix_i_1_25,io_matrix_i_1_24}; // @[RA_Mul.scala 702:21:@3985.4]
  assign _T_1725 = {io_matrix_i_1_27,io_matrix_i_1_26}; // @[RA_Mul.scala 702:21:@3986.4]
  assign _T_1726 = {_T_1725,_T_1724}; // @[RA_Mul.scala 702:21:@3987.4]
  assign _T_1727 = {io_matrix_i_1_29,1'h0}; // @[RA_Mul.scala 702:21:@3988.4]
  assign _T_1728 = {io_matrix_i_1_31,1'h0}; // @[RA_Mul.scala 702:21:@3989.4]
  assign _T_1729 = {_T_1728,_T_1727}; // @[RA_Mul.scala 702:21:@3990.4]
  assign _T_1730 = {_T_1729,_T_1726}; // @[RA_Mul.scala 702:21:@3991.4]
  assign _T_1731 = {_T_1730,_T_1723}; // @[RA_Mul.scala 702:21:@3992.4]
  assign _T_1732 = {_T_1731,_T_1716}; // @[RA_Mul.scala 702:21:@3993.4]
  assign io_matrix_o_0_0 = tmp_0[0]; // @[RA_Mul.scala 705:7:@4029.4]
  assign io_matrix_o_0_1 = tmp_0[1]; // @[RA_Mul.scala 705:7:@4030.4]
  assign io_matrix_o_0_2 = tmp_0[2]; // @[RA_Mul.scala 705:7:@4031.4]
  assign io_matrix_o_0_3 = tmp_0[3]; // @[RA_Mul.scala 705:7:@4032.4]
  assign io_matrix_o_0_4 = tmp_0[4]; // @[RA_Mul.scala 705:7:@4033.4]
  assign io_matrix_o_0_5 = tmp_0[5]; // @[RA_Mul.scala 705:7:@4034.4]
  assign io_matrix_o_0_6 = tmp_0[6]; // @[RA_Mul.scala 705:7:@4035.4]
  assign io_matrix_o_0_7 = tmp_0[7]; // @[RA_Mul.scala 705:7:@4036.4]
  assign io_matrix_o_0_8 = tmp_0[8]; // @[RA_Mul.scala 705:7:@4037.4]
  assign io_matrix_o_0_9 = tmp_0[9]; // @[RA_Mul.scala 705:7:@4038.4]
  assign io_matrix_o_0_10 = tmp_0[10]; // @[RA_Mul.scala 705:7:@4039.4]
  assign io_matrix_o_0_11 = tmp_0[11]; // @[RA_Mul.scala 705:7:@4040.4]
  assign io_matrix_o_0_12 = tmp_0[12]; // @[RA_Mul.scala 705:7:@4041.4]
  assign io_matrix_o_0_13 = tmp_0[13]; // @[RA_Mul.scala 705:7:@4042.4]
  assign io_matrix_o_0_14 = tmp_0[14]; // @[RA_Mul.scala 705:7:@4043.4]
  assign io_matrix_o_0_15 = tmp_0[15]; // @[RA_Mul.scala 705:7:@4044.4]
  assign io_matrix_o_0_16 = tmp_0[16]; // @[RA_Mul.scala 705:7:@4045.4]
  assign io_matrix_o_0_17 = tmp_0[17]; // @[RA_Mul.scala 705:7:@4046.4]
  assign io_matrix_o_0_18 = tmp_0[18]; // @[RA_Mul.scala 705:7:@4047.4]
  assign io_matrix_o_0_19 = tmp_0[19]; // @[RA_Mul.scala 705:7:@4048.4]
  assign io_matrix_o_0_20 = tmp_0[20]; // @[RA_Mul.scala 705:7:@4049.4]
  assign io_matrix_o_0_21 = tmp_0[21]; // @[RA_Mul.scala 705:7:@4050.4]
  assign io_matrix_o_0_22 = tmp_0[22]; // @[RA_Mul.scala 705:7:@4051.4]
  assign io_matrix_o_0_23 = tmp_0[23]; // @[RA_Mul.scala 705:7:@4052.4]
  assign io_matrix_o_0_24 = tmp_0[24]; // @[RA_Mul.scala 705:7:@4053.4]
  assign io_matrix_o_0_25 = tmp_0[25]; // @[RA_Mul.scala 705:7:@4054.4]
  assign io_matrix_o_0_26 = tmp_0[26]; // @[RA_Mul.scala 705:7:@4055.4]
  assign io_matrix_o_0_27 = tmp_0[27]; // @[RA_Mul.scala 705:7:@4056.4]
  assign io_matrix_o_0_28 = tmp_0[28]; // @[RA_Mul.scala 705:7:@4057.4]
  assign io_matrix_o_0_29 = tmp_0[29]; // @[RA_Mul.scala 705:7:@4058.4]
  assign io_matrix_o_0_30 = tmp_0[30]; // @[RA_Mul.scala 705:7:@4059.4]
  assign io_matrix_o_0_31 = tmp_0[31]; // @[RA_Mul.scala 705:7:@4060.4]
  assign io_matrix_o_1_0 = tmp_1[0]; // @[RA_Mul.scala 705:7:@4093.4]
  assign io_matrix_o_1_1 = tmp_1[1]; // @[RA_Mul.scala 705:7:@4094.4]
  assign io_matrix_o_1_2 = tmp_1[2]; // @[RA_Mul.scala 705:7:@4095.4]
  assign io_matrix_o_1_3 = tmp_1[3]; // @[RA_Mul.scala 705:7:@4096.4]
  assign io_matrix_o_1_4 = tmp_1[4]; // @[RA_Mul.scala 705:7:@4097.4]
  assign io_matrix_o_1_5 = tmp_1[5]; // @[RA_Mul.scala 705:7:@4098.4]
  assign io_matrix_o_1_6 = tmp_1[6]; // @[RA_Mul.scala 705:7:@4099.4]
  assign io_matrix_o_1_7 = tmp_1[7]; // @[RA_Mul.scala 705:7:@4100.4]
  assign io_matrix_o_1_8 = tmp_1[8]; // @[RA_Mul.scala 705:7:@4101.4]
  assign io_matrix_o_1_9 = tmp_1[9]; // @[RA_Mul.scala 705:7:@4102.4]
  assign io_matrix_o_1_10 = tmp_1[10]; // @[RA_Mul.scala 705:7:@4103.4]
  assign io_matrix_o_1_11 = tmp_1[11]; // @[RA_Mul.scala 705:7:@4104.4]
  assign io_matrix_o_1_12 = tmp_1[12]; // @[RA_Mul.scala 705:7:@4105.4]
  assign io_matrix_o_1_13 = tmp_1[13]; // @[RA_Mul.scala 705:7:@4106.4]
  assign io_matrix_o_1_14 = tmp_1[14]; // @[RA_Mul.scala 705:7:@4107.4]
  assign io_matrix_o_1_15 = tmp_1[15]; // @[RA_Mul.scala 705:7:@4108.4]
  assign io_matrix_o_1_16 = tmp_1[16]; // @[RA_Mul.scala 705:7:@4109.4]
  assign io_matrix_o_1_17 = tmp_1[17]; // @[RA_Mul.scala 705:7:@4110.4]
  assign io_matrix_o_1_18 = tmp_1[18]; // @[RA_Mul.scala 705:7:@4111.4]
  assign io_matrix_o_1_19 = tmp_1[19]; // @[RA_Mul.scala 705:7:@4112.4]
  assign io_matrix_o_1_20 = tmp_1[20]; // @[RA_Mul.scala 705:7:@4113.4]
  assign io_matrix_o_1_21 = tmp_1[21]; // @[RA_Mul.scala 705:7:@4114.4]
  assign io_matrix_o_1_22 = tmp_1[22]; // @[RA_Mul.scala 705:7:@4115.4]
  assign io_matrix_o_1_23 = tmp_1[23]; // @[RA_Mul.scala 705:7:@4116.4]
  assign io_matrix_o_1_24 = tmp_1[24]; // @[RA_Mul.scala 705:7:@4117.4]
  assign io_matrix_o_1_25 = tmp_1[25]; // @[RA_Mul.scala 705:7:@4118.4]
  assign io_matrix_o_1_26 = tmp_1[26]; // @[RA_Mul.scala 705:7:@4119.4]
  assign io_matrix_o_1_27 = tmp_1[27]; // @[RA_Mul.scala 705:7:@4120.4]
  assign io_matrix_o_1_28 = tmp_1[28]; // @[RA_Mul.scala 705:7:@4121.4]
  assign io_matrix_o_1_29 = tmp_1[29]; // @[RA_Mul.scala 705:7:@4122.4]
  assign io_matrix_o_1_30 = tmp_1[30]; // @[RA_Mul.scala 705:7:@4123.4]
  assign io_matrix_o_1_31 = tmp_1[31]; // @[RA_Mul.scala 705:7:@4124.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tmp_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tmp_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      tmp_0 <= 32'h0;
    end else begin
      tmp_0 <= _T_1698;
    end
    if (reset) begin
      tmp_1 <= 32'h0;
    end else begin
      tmp_1 <= _T_1732;
    end
  end
endmodule
module TailAdder( // @[:@4126.2]
  output [31:0] io_S, // @[:@4129.4]
  input  [31:0] io_B, // @[:@4129.4]
  input  [31:0] io_A // @[:@4129.4]
);
  wire [32:0] _T_11; // @[RA_Mul.scala 612:16:@4131.4]
  assign _T_11 = io_A + io_B; // @[RA_Mul.scala 612:16:@4131.4]
  assign io_S = _T_11[31:0]; // @[RA_Mul.scala 612:8:@4133.4]
endmodule
module PPLRegs3( // @[:@4135.2]
  input         clock, // @[:@4136.4]
  input         reset, // @[:@4137.4]
  output [31:0] io_S_o, // @[:@4138.4]
  input  [31:0] io_S_i // @[:@4138.4]
);
  reg [31:0] _T_11; // @[RA_Mul.scala 724:20:@4140.4]
  reg [31:0] _RAND_0;
  assign io_S_o = _T_11; // @[RA_Mul.scala 724:10:@4142.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_11 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_11 <= 32'h0;
    end else begin
      _T_11 <= io_S_i;
    end
  end
endmodule
module RA_Mul_ppl( // @[:@4144.2]
  input         clock, // @[:@4145.4]
  input         reset, // @[:@4146.4]
  output [31:0] io_P, // @[:@4147.4]
  input  [15:0] io_B, // @[:@4147.4]
  input  [15:0] io_A // @[:@4147.4]
);
  wire [2:0] BoothEncoder_radix4_io_eB_0; // @[RA_Mul.scala 105:21:@4164.4]
  wire [2:0] BoothEncoder_radix4_io_eB_1; // @[RA_Mul.scala 105:21:@4164.4]
  wire [2:0] BoothEncoder_radix4_io_eB_2; // @[RA_Mul.scala 105:21:@4164.4]
  wire [2:0] BoothEncoder_radix4_io_eB_3; // @[RA_Mul.scala 105:21:@4164.4]
  wire [2:0] BoothEncoder_radix4_io_eB_4; // @[RA_Mul.scala 105:21:@4164.4]
  wire [2:0] BoothEncoder_radix4_io_eB_5; // @[RA_Mul.scala 105:21:@4164.4]
  wire [2:0] BoothEncoder_radix4_io_eB_6; // @[RA_Mul.scala 105:21:@4164.4]
  wire [2:0] BoothEncoder_radix4_io_eB_7; // @[RA_Mul.scala 105:21:@4164.4]
  wire [15:0] BoothEncoder_radix4_io_B; // @[RA_Mul.scala 105:21:@4164.4]
  wire [15:0] PPGen_io_PP_0; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_PP_1; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_PP_2; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_PP_3; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_PP_4; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_PP_5; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_PP_6; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_PP_7; // @[RA_Mul.scala 159:21:@4176.4]
  wire [7:0] PPGen_io_SC; // @[RA_Mul.scala 159:21:@4176.4]
  wire [7:0] PPGen_io_S; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_0; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_1; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_2; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_3; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_4; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_5; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_6; // @[RA_Mul.scala 159:21:@4176.4]
  wire [2:0] PPGen_io_eB_7; // @[RA_Mul.scala 159:21:@4176.4]
  wire [15:0] PPGen_io_A; // @[RA_Mul.scala 159:21:@4176.4]
  wire  PPLRegs1_clock; // @[RA_Mul.scala 679:21:@4199.4]
  wire  PPLRegs1_reset; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_0; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_1; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_2; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_3; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_4; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_5; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_6; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_i_7; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_0; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_1; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_2; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_3; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_4; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_5; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_6; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_PP_o_7; // @[RA_Mul.scala 679:21:@4199.4]
  wire [15:0] PPLRegs1_io_SS_o; // @[RA_Mul.scala 679:21:@4199.4]
  wire [7:0] PPLRegs1_io_SC_i; // @[RA_Mul.scala 679:21:@4199.4]
  wire [7:0] PPLRegs1_io_SC_o; // @[RA_Mul.scala 679:21:@4199.4]
  wire [7:0] PPLRegs1_io_S_i; // @[RA_Mul.scala 679:21:@4199.4]
  wire [7:0] PPLRegs1_io_S_o; // @[RA_Mul.scala 679:21:@4199.4]
  wire  Reduction_1_io_matrix_0_0; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_1; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_2; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_3; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_4; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_5; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_6; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_7; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_8; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_9; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_10; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_11; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_12; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_13; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_14; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_15; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_16; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_17; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_18; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_19; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_20; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_21; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_22; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_23; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_24; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_25; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_26; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_27; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_28; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_29; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_30; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_0_31; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_1; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_3; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_4; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_5; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_6; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_7; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_8; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_9; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_10; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_11; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_12; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_13; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_14; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_15; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_16; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_17; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_18; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_19; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_20; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_21; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_22; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_23; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_24; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_25; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_26; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_27; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_28; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_29; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_1_30; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_3; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_6; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_7; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_8; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_9; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_10; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_11; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_12; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_13; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_14; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_15; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_16; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_17; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_18; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_19; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_20; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_21; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_22; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_23; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_24; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_25; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_26; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_2_29; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_6; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_9; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_10; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_11; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_12; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_13; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_14; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_15; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_16; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_17; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_18; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_19; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_20; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_21; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_22; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_23; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_3_24; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_9; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_12; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_13; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_14; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_15; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_16; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_17; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_18; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_19; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_20; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_4_23; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_5_12; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_5_15; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_5_16; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_5_17; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_5_18; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_1_io_matrix_5_19; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_0; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_1; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_2; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_3; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_4; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_5; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_6; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_PP_7; // @[RA_Mul.scala 320:21:@4224.4]
  wire [15:0] Reduction_1_io_SS; // @[RA_Mul.scala 320:21:@4224.4]
  wire [7:0] Reduction_1_io_SC; // @[RA_Mul.scala 320:21:@4224.4]
  wire [7:0] Reduction_1_io_S; // @[RA_Mul.scala 320:21:@4224.4]
  wire  Reduction_2_io_matrix_o_0_0; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_1; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_2; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_3; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_4; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_5; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_6; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_7; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_8; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_10; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_11; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_22; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_24; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_25; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_26; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_27; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_28; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_29; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_30; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_0_31; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_2; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_4; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_5; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_6; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_7; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_8; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_10; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_11; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_22; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_24; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_25; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_26; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_27; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_28; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_1_30; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_4; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_10; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_11; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_22; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_24; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_27; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_2_30; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_o_3_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_0; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_1; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_2; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_3; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_4; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_5; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_6; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_7; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_8; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_10; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_11; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_22; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_24; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_25; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_26; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_27; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_28; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_29; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_30; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_0_31; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_1; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_3; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_4; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_5; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_6; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_7; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_8; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_10; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_11; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_22; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_24; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_25; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_26; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_27; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_28; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_29; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_1_30; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_3; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_6; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_7; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_8; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_10; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_11; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_22; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_24; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_25; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_26; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_2_29; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_6; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_10; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_11; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_21; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_22; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_3_24; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_9; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_13; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_14; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_20; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_4_23; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_5_12; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_5_15; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_5_16; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_5_17; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_5_18; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_2_io_matrix_i_5_19; // @[RA_Mul.scala 444:21:@4430.4]
  wire  Reduction_3_io_matrix_o_0_0; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_1; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_2; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_3; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_4; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_5; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_6; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_7; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_8; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_9; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_10; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_11; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_12; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_13; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_14; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_15; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_16; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_17; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_18; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_19; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_20; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_21; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_22; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_23; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_24; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_25; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_26; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_27; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_28; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_29; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_30; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_0_31; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_3; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_5; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_6; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_7; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_8; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_9; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_10; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_11; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_12; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_13; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_14; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_15; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_16; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_17; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_18; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_19; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_20; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_21; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_22; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_23; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_24; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_25; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_26; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_28; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_1_31; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_5; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_13; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_14; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_15; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_16; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_17; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_18; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_19; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_20; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_21; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_23; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_25; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_o_2_28; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_0; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_1; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_2; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_3; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_4; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_5; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_6; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_7; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_8; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_9; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_10; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_11; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_12; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_13; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_14; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_15; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_16; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_17; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_18; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_19; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_20; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_21; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_22; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_23; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_24; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_25; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_26; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_27; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_28; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_29; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_30; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_0_31; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_2; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_4; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_5; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_6; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_7; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_8; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_9; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_10; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_11; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_12; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_13; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_14; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_15; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_16; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_17; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_18; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_19; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_20; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_21; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_22; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_23; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_24; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_25; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_26; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_27; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_28; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_1_30; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_4; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_9; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_10; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_11; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_12; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_13; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_14; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_15; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_16; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_17; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_18; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_19; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_20; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_21; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_22; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_23; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_24; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_27; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_2_30; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_9; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_13; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_14; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_15; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_16; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_17; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_18; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_19; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_20; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_21; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_3_io_matrix_i_3_23; // @[RA_Mul.scala 535:21:@4753.4]
  wire  Reduction_4_io_matrix_o_0_0; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_1; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_2; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_3; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_4; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_5; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_6; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_7; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_8; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_9; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_10; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_11; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_12; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_13; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_14; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_15; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_16; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_17; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_18; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_19; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_20; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_21; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_22; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_23; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_24; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_25; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_26; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_27; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_28; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_29; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_30; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_0_31; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_4; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_6; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_7; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_8; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_9; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_10; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_11; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_12; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_13; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_14; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_15; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_16; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_17; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_18; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_19; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_20; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_21; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_22; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_23; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_24; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_25; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_26; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_27; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_29; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_o_1_31; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_0; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_1; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_2; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_3; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_4; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_5; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_6; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_7; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_8; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_9; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_10; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_11; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_12; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_13; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_14; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_15; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_16; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_17; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_18; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_19; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_20; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_21; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_22; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_23; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_24; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_25; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_26; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_27; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_28; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_29; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_30; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_0_31; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_3; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_5; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_6; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_7; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_8; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_9; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_10; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_11; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_12; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_13; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_14; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_15; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_16; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_17; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_18; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_19; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_20; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_21; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_22; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_23; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_24; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_25; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_26; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_28; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_1_31; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_5; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_13; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_14; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_15; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_16; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_17; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_18; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_19; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_20; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_21; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_23; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_25; // @[RA_Mul.scala 598:21:@4980.4]
  wire  Reduction_4_io_matrix_i_2_28; // @[RA_Mul.scala 598:21:@4980.4]
  wire  PPLRegs2_clock; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_reset; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_0; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_1; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_2; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_3; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_4; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_5; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_6; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_7; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_8; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_9; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_10; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_11; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_12; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_13; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_14; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_15; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_16; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_17; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_18; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_19; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_20; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_21; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_22; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_23; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_24; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_25; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_26; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_27; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_28; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_29; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_30; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_0_31; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_0; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_1; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_2; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_3; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_4; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_5; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_6; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_7; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_8; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_9; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_10; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_11; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_12; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_13; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_14; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_15; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_16; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_17; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_18; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_19; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_20; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_21; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_22; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_23; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_24; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_25; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_26; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_27; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_28; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_29; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_30; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_o_1_31; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_0; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_1; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_2; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_3; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_4; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_5; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_6; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_7; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_8; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_9; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_10; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_11; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_12; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_13; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_14; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_15; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_16; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_17; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_18; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_19; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_20; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_21; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_22; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_23; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_24; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_25; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_26; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_27; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_28; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_29; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_30; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_0_31; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_4; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_6; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_7; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_8; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_9; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_10; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_11; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_12; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_13; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_14; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_15; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_16; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_17; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_18; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_19; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_20; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_21; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_22; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_23; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_24; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_25; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_26; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_27; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_29; // @[RA_Mul.scala 711:21:@5143.4]
  wire  PPLRegs2_io_matrix_i_1_31; // @[RA_Mul.scala 711:21:@5143.4]
  wire [31:0] TailAdder_io_S; // @[RA_Mul.scala 617:21:@5336.4]
  wire [31:0] TailAdder_io_B; // @[RA_Mul.scala 617:21:@5336.4]
  wire [31:0] TailAdder_io_A; // @[RA_Mul.scala 617:21:@5336.4]
  wire  PPLRegs3_clock; // @[RA_Mul.scala 729:21:@5342.4]
  wire  PPLRegs3_reset; // @[RA_Mul.scala 729:21:@5342.4]
  wire [31:0] PPLRegs3_io_S_o; // @[RA_Mul.scala 729:21:@5342.4]
  wire [31:0] PPLRegs3_io_S_i; // @[RA_Mul.scala 729:21:@5342.4]
  wire  matrix_o4_o_0_1; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5147.4]
  wire  matrix_o4_o_0_0; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5146.4]
  wire [1:0] _T_3079; // @[RA_Mul.scala 769:28:@5274.4]
  wire  matrix_o4_o_0_3; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5149.4]
  wire  matrix_o4_o_0_2; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5148.4]
  wire [1:0] _T_3080; // @[RA_Mul.scala 769:28:@5275.4]
  wire [3:0] _T_3081; // @[RA_Mul.scala 769:28:@5276.4]
  wire  matrix_o4_o_0_5; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5151.4]
  wire  matrix_o4_o_0_4; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5150.4]
  wire [1:0] _T_3082; // @[RA_Mul.scala 769:28:@5277.4]
  wire  matrix_o4_o_0_7; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5153.4]
  wire  matrix_o4_o_0_6; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5152.4]
  wire [1:0] _T_3083; // @[RA_Mul.scala 769:28:@5278.4]
  wire [3:0] _T_3084; // @[RA_Mul.scala 769:28:@5279.4]
  wire [7:0] _T_3085; // @[RA_Mul.scala 769:28:@5280.4]
  wire  matrix_o4_o_0_9; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5155.4]
  wire  matrix_o4_o_0_8; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5154.4]
  wire [1:0] _T_3086; // @[RA_Mul.scala 769:28:@5281.4]
  wire  matrix_o4_o_0_11; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5157.4]
  wire  matrix_o4_o_0_10; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5156.4]
  wire [1:0] _T_3087; // @[RA_Mul.scala 769:28:@5282.4]
  wire [3:0] _T_3088; // @[RA_Mul.scala 769:28:@5283.4]
  wire  matrix_o4_o_0_13; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5159.4]
  wire  matrix_o4_o_0_12; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5158.4]
  wire [1:0] _T_3089; // @[RA_Mul.scala 769:28:@5284.4]
  wire  matrix_o4_o_0_15; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5161.4]
  wire  matrix_o4_o_0_14; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5160.4]
  wire [1:0] _T_3090; // @[RA_Mul.scala 769:28:@5285.4]
  wire [3:0] _T_3091; // @[RA_Mul.scala 769:28:@5286.4]
  wire [7:0] _T_3092; // @[RA_Mul.scala 769:28:@5287.4]
  wire [15:0] _T_3093; // @[RA_Mul.scala 769:28:@5288.4]
  wire  matrix_o4_o_0_17; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5163.4]
  wire  matrix_o4_o_0_16; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5162.4]
  wire [1:0] _T_3094; // @[RA_Mul.scala 769:28:@5289.4]
  wire  matrix_o4_o_0_19; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5165.4]
  wire  matrix_o4_o_0_18; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5164.4]
  wire [1:0] _T_3095; // @[RA_Mul.scala 769:28:@5290.4]
  wire [3:0] _T_3096; // @[RA_Mul.scala 769:28:@5291.4]
  wire  matrix_o4_o_0_21; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5167.4]
  wire  matrix_o4_o_0_20; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5166.4]
  wire [1:0] _T_3097; // @[RA_Mul.scala 769:28:@5292.4]
  wire  matrix_o4_o_0_23; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5169.4]
  wire  matrix_o4_o_0_22; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5168.4]
  wire [1:0] _T_3098; // @[RA_Mul.scala 769:28:@5293.4]
  wire [3:0] _T_3099; // @[RA_Mul.scala 769:28:@5294.4]
  wire [7:0] _T_3100; // @[RA_Mul.scala 769:28:@5295.4]
  wire  matrix_o4_o_0_25; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5171.4]
  wire  matrix_o4_o_0_24; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5170.4]
  wire [1:0] _T_3101; // @[RA_Mul.scala 769:28:@5296.4]
  wire  matrix_o4_o_0_27; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5173.4]
  wire  matrix_o4_o_0_26; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5172.4]
  wire [1:0] _T_3102; // @[RA_Mul.scala 769:28:@5297.4]
  wire [3:0] _T_3103; // @[RA_Mul.scala 769:28:@5298.4]
  wire  matrix_o4_o_0_29; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5175.4]
  wire  matrix_o4_o_0_28; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5174.4]
  wire [1:0] _T_3104; // @[RA_Mul.scala 769:28:@5299.4]
  wire  matrix_o4_o_0_31; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5177.4]
  wire  matrix_o4_o_0_30; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5176.4]
  wire [1:0] _T_3105; // @[RA_Mul.scala 769:28:@5300.4]
  wire [3:0] _T_3106; // @[RA_Mul.scala 769:28:@5301.4]
  wire [7:0] _T_3107; // @[RA_Mul.scala 769:28:@5302.4]
  wire [15:0] _T_3108; // @[RA_Mul.scala 769:28:@5303.4]
  wire  matrix_o4_o_1_1; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5179.4]
  wire  matrix_o4_o_1_0; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5178.4]
  wire [1:0] _T_3110; // @[RA_Mul.scala 769:51:@5305.4]
  wire  matrix_o4_o_1_3; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5181.4]
  wire  matrix_o4_o_1_2; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5180.4]
  wire [1:0] _T_3111; // @[RA_Mul.scala 769:51:@5306.4]
  wire [3:0] _T_3112; // @[RA_Mul.scala 769:51:@5307.4]
  wire  matrix_o4_o_1_5; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5183.4]
  wire  matrix_o4_o_1_4; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5182.4]
  wire [1:0] _T_3113; // @[RA_Mul.scala 769:51:@5308.4]
  wire  matrix_o4_o_1_7; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5185.4]
  wire  matrix_o4_o_1_6; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5184.4]
  wire [1:0] _T_3114; // @[RA_Mul.scala 769:51:@5309.4]
  wire [3:0] _T_3115; // @[RA_Mul.scala 769:51:@5310.4]
  wire [7:0] _T_3116; // @[RA_Mul.scala 769:51:@5311.4]
  wire  matrix_o4_o_1_9; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5187.4]
  wire  matrix_o4_o_1_8; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5186.4]
  wire [1:0] _T_3117; // @[RA_Mul.scala 769:51:@5312.4]
  wire  matrix_o4_o_1_11; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5189.4]
  wire  matrix_o4_o_1_10; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5188.4]
  wire [1:0] _T_3118; // @[RA_Mul.scala 769:51:@5313.4]
  wire [3:0] _T_3119; // @[RA_Mul.scala 769:51:@5314.4]
  wire  matrix_o4_o_1_13; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5191.4]
  wire  matrix_o4_o_1_12; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5190.4]
  wire [1:0] _T_3120; // @[RA_Mul.scala 769:51:@5315.4]
  wire  matrix_o4_o_1_15; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5193.4]
  wire  matrix_o4_o_1_14; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5192.4]
  wire [1:0] _T_3121; // @[RA_Mul.scala 769:51:@5316.4]
  wire [3:0] _T_3122; // @[RA_Mul.scala 769:51:@5317.4]
  wire [7:0] _T_3123; // @[RA_Mul.scala 769:51:@5318.4]
  wire [15:0] _T_3124; // @[RA_Mul.scala 769:51:@5319.4]
  wire  matrix_o4_o_1_17; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5195.4]
  wire  matrix_o4_o_1_16; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5194.4]
  wire [1:0] _T_3125; // @[RA_Mul.scala 769:51:@5320.4]
  wire  matrix_o4_o_1_19; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5197.4]
  wire  matrix_o4_o_1_18; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5196.4]
  wire [1:0] _T_3126; // @[RA_Mul.scala 769:51:@5321.4]
  wire [3:0] _T_3127; // @[RA_Mul.scala 769:51:@5322.4]
  wire  matrix_o4_o_1_21; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5199.4]
  wire  matrix_o4_o_1_20; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5198.4]
  wire [1:0] _T_3128; // @[RA_Mul.scala 769:51:@5323.4]
  wire  matrix_o4_o_1_23; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5201.4]
  wire  matrix_o4_o_1_22; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5200.4]
  wire [1:0] _T_3129; // @[RA_Mul.scala 769:51:@5324.4]
  wire [3:0] _T_3130; // @[RA_Mul.scala 769:51:@5325.4]
  wire [7:0] _T_3131; // @[RA_Mul.scala 769:51:@5326.4]
  wire  matrix_o4_o_1_25; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5203.4]
  wire  matrix_o4_o_1_24; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5202.4]
  wire [1:0] _T_3132; // @[RA_Mul.scala 769:51:@5327.4]
  wire  matrix_o4_o_1_27; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5205.4]
  wire  matrix_o4_o_1_26; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5204.4]
  wire [1:0] _T_3133; // @[RA_Mul.scala 769:51:@5328.4]
  wire [3:0] _T_3134; // @[RA_Mul.scala 769:51:@5329.4]
  wire  matrix_o4_o_1_29; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5207.4]
  wire  matrix_o4_o_1_28; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5206.4]
  wire [1:0] _T_3135; // @[RA_Mul.scala 769:51:@5330.4]
  wire  matrix_o4_o_1_31; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5209.4]
  wire  matrix_o4_o_1_30; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5208.4]
  wire [1:0] _T_3136; // @[RA_Mul.scala 769:51:@5331.4]
  wire [3:0] _T_3137; // @[RA_Mul.scala 769:51:@5332.4]
  wire [7:0] _T_3138; // @[RA_Mul.scala 769:51:@5333.4]
  wire [15:0] _T_3139; // @[RA_Mul.scala 769:51:@5334.4]
  BoothEncoder_radix4 BoothEncoder_radix4 ( // @[RA_Mul.scala 105:21:@4164.4]
    .io_eB_0(BoothEncoder_radix4_io_eB_0),
    .io_eB_1(BoothEncoder_radix4_io_eB_1),
    .io_eB_2(BoothEncoder_radix4_io_eB_2),
    .io_eB_3(BoothEncoder_radix4_io_eB_3),
    .io_eB_4(BoothEncoder_radix4_io_eB_4),
    .io_eB_5(BoothEncoder_radix4_io_eB_5),
    .io_eB_6(BoothEncoder_radix4_io_eB_6),
    .io_eB_7(BoothEncoder_radix4_io_eB_7),
    .io_B(BoothEncoder_radix4_io_B)
  );
  PPGen PPGen ( // @[RA_Mul.scala 159:21:@4176.4]
    .io_PP_0(PPGen_io_PP_0),
    .io_PP_1(PPGen_io_PP_1),
    .io_PP_2(PPGen_io_PP_2),
    .io_PP_3(PPGen_io_PP_3),
    .io_PP_4(PPGen_io_PP_4),
    .io_PP_5(PPGen_io_PP_5),
    .io_PP_6(PPGen_io_PP_6),
    .io_PP_7(PPGen_io_PP_7),
    .io_SC(PPGen_io_SC),
    .io_S(PPGen_io_S),
    .io_eB_0(PPGen_io_eB_0),
    .io_eB_1(PPGen_io_eB_1),
    .io_eB_2(PPGen_io_eB_2),
    .io_eB_3(PPGen_io_eB_3),
    .io_eB_4(PPGen_io_eB_4),
    .io_eB_5(PPGen_io_eB_5),
    .io_eB_6(PPGen_io_eB_6),
    .io_eB_7(PPGen_io_eB_7),
    .io_A(PPGen_io_A)
  );
  PPLRegs1 PPLRegs1 ( // @[RA_Mul.scala 679:21:@4199.4]
    .clock(PPLRegs1_clock),
    .reset(PPLRegs1_reset),
    .io_PP_i_0(PPLRegs1_io_PP_i_0),
    .io_PP_i_1(PPLRegs1_io_PP_i_1),
    .io_PP_i_2(PPLRegs1_io_PP_i_2),
    .io_PP_i_3(PPLRegs1_io_PP_i_3),
    .io_PP_i_4(PPLRegs1_io_PP_i_4),
    .io_PP_i_5(PPLRegs1_io_PP_i_5),
    .io_PP_i_6(PPLRegs1_io_PP_i_6),
    .io_PP_i_7(PPLRegs1_io_PP_i_7),
    .io_PP_o_0(PPLRegs1_io_PP_o_0),
    .io_PP_o_1(PPLRegs1_io_PP_o_1),
    .io_PP_o_2(PPLRegs1_io_PP_o_2),
    .io_PP_o_3(PPLRegs1_io_PP_o_3),
    .io_PP_o_4(PPLRegs1_io_PP_o_4),
    .io_PP_o_5(PPLRegs1_io_PP_o_5),
    .io_PP_o_6(PPLRegs1_io_PP_o_6),
    .io_PP_o_7(PPLRegs1_io_PP_o_7),
    .io_SS_o(PPLRegs1_io_SS_o),
    .io_SC_i(PPLRegs1_io_SC_i),
    .io_SC_o(PPLRegs1_io_SC_o),
    .io_S_i(PPLRegs1_io_S_i),
    .io_S_o(PPLRegs1_io_S_o)
  );
  Reduction_1 Reduction_1 ( // @[RA_Mul.scala 320:21:@4224.4]
    .io_matrix_0_0(Reduction_1_io_matrix_0_0),
    .io_matrix_0_1(Reduction_1_io_matrix_0_1),
    .io_matrix_0_2(Reduction_1_io_matrix_0_2),
    .io_matrix_0_3(Reduction_1_io_matrix_0_3),
    .io_matrix_0_4(Reduction_1_io_matrix_0_4),
    .io_matrix_0_5(Reduction_1_io_matrix_0_5),
    .io_matrix_0_6(Reduction_1_io_matrix_0_6),
    .io_matrix_0_7(Reduction_1_io_matrix_0_7),
    .io_matrix_0_8(Reduction_1_io_matrix_0_8),
    .io_matrix_0_9(Reduction_1_io_matrix_0_9),
    .io_matrix_0_10(Reduction_1_io_matrix_0_10),
    .io_matrix_0_11(Reduction_1_io_matrix_0_11),
    .io_matrix_0_12(Reduction_1_io_matrix_0_12),
    .io_matrix_0_13(Reduction_1_io_matrix_0_13),
    .io_matrix_0_14(Reduction_1_io_matrix_0_14),
    .io_matrix_0_15(Reduction_1_io_matrix_0_15),
    .io_matrix_0_16(Reduction_1_io_matrix_0_16),
    .io_matrix_0_17(Reduction_1_io_matrix_0_17),
    .io_matrix_0_18(Reduction_1_io_matrix_0_18),
    .io_matrix_0_19(Reduction_1_io_matrix_0_19),
    .io_matrix_0_20(Reduction_1_io_matrix_0_20),
    .io_matrix_0_21(Reduction_1_io_matrix_0_21),
    .io_matrix_0_22(Reduction_1_io_matrix_0_22),
    .io_matrix_0_23(Reduction_1_io_matrix_0_23),
    .io_matrix_0_24(Reduction_1_io_matrix_0_24),
    .io_matrix_0_25(Reduction_1_io_matrix_0_25),
    .io_matrix_0_26(Reduction_1_io_matrix_0_26),
    .io_matrix_0_27(Reduction_1_io_matrix_0_27),
    .io_matrix_0_28(Reduction_1_io_matrix_0_28),
    .io_matrix_0_29(Reduction_1_io_matrix_0_29),
    .io_matrix_0_30(Reduction_1_io_matrix_0_30),
    .io_matrix_0_31(Reduction_1_io_matrix_0_31),
    .io_matrix_1_1(Reduction_1_io_matrix_1_1),
    .io_matrix_1_3(Reduction_1_io_matrix_1_3),
    .io_matrix_1_4(Reduction_1_io_matrix_1_4),
    .io_matrix_1_5(Reduction_1_io_matrix_1_5),
    .io_matrix_1_6(Reduction_1_io_matrix_1_6),
    .io_matrix_1_7(Reduction_1_io_matrix_1_7),
    .io_matrix_1_8(Reduction_1_io_matrix_1_8),
    .io_matrix_1_9(Reduction_1_io_matrix_1_9),
    .io_matrix_1_10(Reduction_1_io_matrix_1_10),
    .io_matrix_1_11(Reduction_1_io_matrix_1_11),
    .io_matrix_1_12(Reduction_1_io_matrix_1_12),
    .io_matrix_1_13(Reduction_1_io_matrix_1_13),
    .io_matrix_1_14(Reduction_1_io_matrix_1_14),
    .io_matrix_1_15(Reduction_1_io_matrix_1_15),
    .io_matrix_1_16(Reduction_1_io_matrix_1_16),
    .io_matrix_1_17(Reduction_1_io_matrix_1_17),
    .io_matrix_1_18(Reduction_1_io_matrix_1_18),
    .io_matrix_1_19(Reduction_1_io_matrix_1_19),
    .io_matrix_1_20(Reduction_1_io_matrix_1_20),
    .io_matrix_1_21(Reduction_1_io_matrix_1_21),
    .io_matrix_1_22(Reduction_1_io_matrix_1_22),
    .io_matrix_1_23(Reduction_1_io_matrix_1_23),
    .io_matrix_1_24(Reduction_1_io_matrix_1_24),
    .io_matrix_1_25(Reduction_1_io_matrix_1_25),
    .io_matrix_1_26(Reduction_1_io_matrix_1_26),
    .io_matrix_1_27(Reduction_1_io_matrix_1_27),
    .io_matrix_1_28(Reduction_1_io_matrix_1_28),
    .io_matrix_1_29(Reduction_1_io_matrix_1_29),
    .io_matrix_1_30(Reduction_1_io_matrix_1_30),
    .io_matrix_2_3(Reduction_1_io_matrix_2_3),
    .io_matrix_2_6(Reduction_1_io_matrix_2_6),
    .io_matrix_2_7(Reduction_1_io_matrix_2_7),
    .io_matrix_2_8(Reduction_1_io_matrix_2_8),
    .io_matrix_2_9(Reduction_1_io_matrix_2_9),
    .io_matrix_2_10(Reduction_1_io_matrix_2_10),
    .io_matrix_2_11(Reduction_1_io_matrix_2_11),
    .io_matrix_2_12(Reduction_1_io_matrix_2_12),
    .io_matrix_2_13(Reduction_1_io_matrix_2_13),
    .io_matrix_2_14(Reduction_1_io_matrix_2_14),
    .io_matrix_2_15(Reduction_1_io_matrix_2_15),
    .io_matrix_2_16(Reduction_1_io_matrix_2_16),
    .io_matrix_2_17(Reduction_1_io_matrix_2_17),
    .io_matrix_2_18(Reduction_1_io_matrix_2_18),
    .io_matrix_2_19(Reduction_1_io_matrix_2_19),
    .io_matrix_2_20(Reduction_1_io_matrix_2_20),
    .io_matrix_2_21(Reduction_1_io_matrix_2_21),
    .io_matrix_2_22(Reduction_1_io_matrix_2_22),
    .io_matrix_2_23(Reduction_1_io_matrix_2_23),
    .io_matrix_2_24(Reduction_1_io_matrix_2_24),
    .io_matrix_2_25(Reduction_1_io_matrix_2_25),
    .io_matrix_2_26(Reduction_1_io_matrix_2_26),
    .io_matrix_2_29(Reduction_1_io_matrix_2_29),
    .io_matrix_3_6(Reduction_1_io_matrix_3_6),
    .io_matrix_3_9(Reduction_1_io_matrix_3_9),
    .io_matrix_3_10(Reduction_1_io_matrix_3_10),
    .io_matrix_3_11(Reduction_1_io_matrix_3_11),
    .io_matrix_3_12(Reduction_1_io_matrix_3_12),
    .io_matrix_3_13(Reduction_1_io_matrix_3_13),
    .io_matrix_3_14(Reduction_1_io_matrix_3_14),
    .io_matrix_3_15(Reduction_1_io_matrix_3_15),
    .io_matrix_3_16(Reduction_1_io_matrix_3_16),
    .io_matrix_3_17(Reduction_1_io_matrix_3_17),
    .io_matrix_3_18(Reduction_1_io_matrix_3_18),
    .io_matrix_3_19(Reduction_1_io_matrix_3_19),
    .io_matrix_3_20(Reduction_1_io_matrix_3_20),
    .io_matrix_3_21(Reduction_1_io_matrix_3_21),
    .io_matrix_3_22(Reduction_1_io_matrix_3_22),
    .io_matrix_3_23(Reduction_1_io_matrix_3_23),
    .io_matrix_3_24(Reduction_1_io_matrix_3_24),
    .io_matrix_4_9(Reduction_1_io_matrix_4_9),
    .io_matrix_4_12(Reduction_1_io_matrix_4_12),
    .io_matrix_4_13(Reduction_1_io_matrix_4_13),
    .io_matrix_4_14(Reduction_1_io_matrix_4_14),
    .io_matrix_4_15(Reduction_1_io_matrix_4_15),
    .io_matrix_4_16(Reduction_1_io_matrix_4_16),
    .io_matrix_4_17(Reduction_1_io_matrix_4_17),
    .io_matrix_4_18(Reduction_1_io_matrix_4_18),
    .io_matrix_4_19(Reduction_1_io_matrix_4_19),
    .io_matrix_4_20(Reduction_1_io_matrix_4_20),
    .io_matrix_4_23(Reduction_1_io_matrix_4_23),
    .io_matrix_5_12(Reduction_1_io_matrix_5_12),
    .io_matrix_5_15(Reduction_1_io_matrix_5_15),
    .io_matrix_5_16(Reduction_1_io_matrix_5_16),
    .io_matrix_5_17(Reduction_1_io_matrix_5_17),
    .io_matrix_5_18(Reduction_1_io_matrix_5_18),
    .io_matrix_5_19(Reduction_1_io_matrix_5_19),
    .io_PP_0(Reduction_1_io_PP_0),
    .io_PP_1(Reduction_1_io_PP_1),
    .io_PP_2(Reduction_1_io_PP_2),
    .io_PP_3(Reduction_1_io_PP_3),
    .io_PP_4(Reduction_1_io_PP_4),
    .io_PP_5(Reduction_1_io_PP_5),
    .io_PP_6(Reduction_1_io_PP_6),
    .io_PP_7(Reduction_1_io_PP_7),
    .io_SS(Reduction_1_io_SS),
    .io_SC(Reduction_1_io_SC),
    .io_S(Reduction_1_io_S)
  );
  Reduction_2 Reduction_2 ( // @[RA_Mul.scala 444:21:@4430.4]
    .io_matrix_o_0_0(Reduction_2_io_matrix_o_0_0),
    .io_matrix_o_0_1(Reduction_2_io_matrix_o_0_1),
    .io_matrix_o_0_2(Reduction_2_io_matrix_o_0_2),
    .io_matrix_o_0_3(Reduction_2_io_matrix_o_0_3),
    .io_matrix_o_0_4(Reduction_2_io_matrix_o_0_4),
    .io_matrix_o_0_5(Reduction_2_io_matrix_o_0_5),
    .io_matrix_o_0_6(Reduction_2_io_matrix_o_0_6),
    .io_matrix_o_0_7(Reduction_2_io_matrix_o_0_7),
    .io_matrix_o_0_8(Reduction_2_io_matrix_o_0_8),
    .io_matrix_o_0_9(Reduction_2_io_matrix_o_0_9),
    .io_matrix_o_0_10(Reduction_2_io_matrix_o_0_10),
    .io_matrix_o_0_11(Reduction_2_io_matrix_o_0_11),
    .io_matrix_o_0_12(Reduction_2_io_matrix_o_0_12),
    .io_matrix_o_0_13(Reduction_2_io_matrix_o_0_13),
    .io_matrix_o_0_14(Reduction_2_io_matrix_o_0_14),
    .io_matrix_o_0_15(Reduction_2_io_matrix_o_0_15),
    .io_matrix_o_0_16(Reduction_2_io_matrix_o_0_16),
    .io_matrix_o_0_17(Reduction_2_io_matrix_o_0_17),
    .io_matrix_o_0_18(Reduction_2_io_matrix_o_0_18),
    .io_matrix_o_0_19(Reduction_2_io_matrix_o_0_19),
    .io_matrix_o_0_20(Reduction_2_io_matrix_o_0_20),
    .io_matrix_o_0_21(Reduction_2_io_matrix_o_0_21),
    .io_matrix_o_0_22(Reduction_2_io_matrix_o_0_22),
    .io_matrix_o_0_23(Reduction_2_io_matrix_o_0_23),
    .io_matrix_o_0_24(Reduction_2_io_matrix_o_0_24),
    .io_matrix_o_0_25(Reduction_2_io_matrix_o_0_25),
    .io_matrix_o_0_26(Reduction_2_io_matrix_o_0_26),
    .io_matrix_o_0_27(Reduction_2_io_matrix_o_0_27),
    .io_matrix_o_0_28(Reduction_2_io_matrix_o_0_28),
    .io_matrix_o_0_29(Reduction_2_io_matrix_o_0_29),
    .io_matrix_o_0_30(Reduction_2_io_matrix_o_0_30),
    .io_matrix_o_0_31(Reduction_2_io_matrix_o_0_31),
    .io_matrix_o_1_2(Reduction_2_io_matrix_o_1_2),
    .io_matrix_o_1_4(Reduction_2_io_matrix_o_1_4),
    .io_matrix_o_1_5(Reduction_2_io_matrix_o_1_5),
    .io_matrix_o_1_6(Reduction_2_io_matrix_o_1_6),
    .io_matrix_o_1_7(Reduction_2_io_matrix_o_1_7),
    .io_matrix_o_1_8(Reduction_2_io_matrix_o_1_8),
    .io_matrix_o_1_9(Reduction_2_io_matrix_o_1_9),
    .io_matrix_o_1_10(Reduction_2_io_matrix_o_1_10),
    .io_matrix_o_1_11(Reduction_2_io_matrix_o_1_11),
    .io_matrix_o_1_12(Reduction_2_io_matrix_o_1_12),
    .io_matrix_o_1_13(Reduction_2_io_matrix_o_1_13),
    .io_matrix_o_1_14(Reduction_2_io_matrix_o_1_14),
    .io_matrix_o_1_15(Reduction_2_io_matrix_o_1_15),
    .io_matrix_o_1_16(Reduction_2_io_matrix_o_1_16),
    .io_matrix_o_1_17(Reduction_2_io_matrix_o_1_17),
    .io_matrix_o_1_18(Reduction_2_io_matrix_o_1_18),
    .io_matrix_o_1_19(Reduction_2_io_matrix_o_1_19),
    .io_matrix_o_1_20(Reduction_2_io_matrix_o_1_20),
    .io_matrix_o_1_21(Reduction_2_io_matrix_o_1_21),
    .io_matrix_o_1_22(Reduction_2_io_matrix_o_1_22),
    .io_matrix_o_1_23(Reduction_2_io_matrix_o_1_23),
    .io_matrix_o_1_24(Reduction_2_io_matrix_o_1_24),
    .io_matrix_o_1_25(Reduction_2_io_matrix_o_1_25),
    .io_matrix_o_1_26(Reduction_2_io_matrix_o_1_26),
    .io_matrix_o_1_27(Reduction_2_io_matrix_o_1_27),
    .io_matrix_o_1_28(Reduction_2_io_matrix_o_1_28),
    .io_matrix_o_1_30(Reduction_2_io_matrix_o_1_30),
    .io_matrix_o_2_4(Reduction_2_io_matrix_o_2_4),
    .io_matrix_o_2_9(Reduction_2_io_matrix_o_2_9),
    .io_matrix_o_2_10(Reduction_2_io_matrix_o_2_10),
    .io_matrix_o_2_11(Reduction_2_io_matrix_o_2_11),
    .io_matrix_o_2_12(Reduction_2_io_matrix_o_2_12),
    .io_matrix_o_2_13(Reduction_2_io_matrix_o_2_13),
    .io_matrix_o_2_14(Reduction_2_io_matrix_o_2_14),
    .io_matrix_o_2_15(Reduction_2_io_matrix_o_2_15),
    .io_matrix_o_2_16(Reduction_2_io_matrix_o_2_16),
    .io_matrix_o_2_17(Reduction_2_io_matrix_o_2_17),
    .io_matrix_o_2_18(Reduction_2_io_matrix_o_2_18),
    .io_matrix_o_2_19(Reduction_2_io_matrix_o_2_19),
    .io_matrix_o_2_20(Reduction_2_io_matrix_o_2_20),
    .io_matrix_o_2_21(Reduction_2_io_matrix_o_2_21),
    .io_matrix_o_2_22(Reduction_2_io_matrix_o_2_22),
    .io_matrix_o_2_23(Reduction_2_io_matrix_o_2_23),
    .io_matrix_o_2_24(Reduction_2_io_matrix_o_2_24),
    .io_matrix_o_2_27(Reduction_2_io_matrix_o_2_27),
    .io_matrix_o_2_30(Reduction_2_io_matrix_o_2_30),
    .io_matrix_o_3_9(Reduction_2_io_matrix_o_3_9),
    .io_matrix_o_3_13(Reduction_2_io_matrix_o_3_13),
    .io_matrix_o_3_14(Reduction_2_io_matrix_o_3_14),
    .io_matrix_o_3_15(Reduction_2_io_matrix_o_3_15),
    .io_matrix_o_3_16(Reduction_2_io_matrix_o_3_16),
    .io_matrix_o_3_17(Reduction_2_io_matrix_o_3_17),
    .io_matrix_o_3_18(Reduction_2_io_matrix_o_3_18),
    .io_matrix_o_3_19(Reduction_2_io_matrix_o_3_19),
    .io_matrix_o_3_20(Reduction_2_io_matrix_o_3_20),
    .io_matrix_o_3_21(Reduction_2_io_matrix_o_3_21),
    .io_matrix_o_3_23(Reduction_2_io_matrix_o_3_23),
    .io_matrix_i_0_0(Reduction_2_io_matrix_i_0_0),
    .io_matrix_i_0_1(Reduction_2_io_matrix_i_0_1),
    .io_matrix_i_0_2(Reduction_2_io_matrix_i_0_2),
    .io_matrix_i_0_3(Reduction_2_io_matrix_i_0_3),
    .io_matrix_i_0_4(Reduction_2_io_matrix_i_0_4),
    .io_matrix_i_0_5(Reduction_2_io_matrix_i_0_5),
    .io_matrix_i_0_6(Reduction_2_io_matrix_i_0_6),
    .io_matrix_i_0_7(Reduction_2_io_matrix_i_0_7),
    .io_matrix_i_0_8(Reduction_2_io_matrix_i_0_8),
    .io_matrix_i_0_9(Reduction_2_io_matrix_i_0_9),
    .io_matrix_i_0_10(Reduction_2_io_matrix_i_0_10),
    .io_matrix_i_0_11(Reduction_2_io_matrix_i_0_11),
    .io_matrix_i_0_12(Reduction_2_io_matrix_i_0_12),
    .io_matrix_i_0_13(Reduction_2_io_matrix_i_0_13),
    .io_matrix_i_0_14(Reduction_2_io_matrix_i_0_14),
    .io_matrix_i_0_15(Reduction_2_io_matrix_i_0_15),
    .io_matrix_i_0_16(Reduction_2_io_matrix_i_0_16),
    .io_matrix_i_0_17(Reduction_2_io_matrix_i_0_17),
    .io_matrix_i_0_18(Reduction_2_io_matrix_i_0_18),
    .io_matrix_i_0_19(Reduction_2_io_matrix_i_0_19),
    .io_matrix_i_0_20(Reduction_2_io_matrix_i_0_20),
    .io_matrix_i_0_21(Reduction_2_io_matrix_i_0_21),
    .io_matrix_i_0_22(Reduction_2_io_matrix_i_0_22),
    .io_matrix_i_0_23(Reduction_2_io_matrix_i_0_23),
    .io_matrix_i_0_24(Reduction_2_io_matrix_i_0_24),
    .io_matrix_i_0_25(Reduction_2_io_matrix_i_0_25),
    .io_matrix_i_0_26(Reduction_2_io_matrix_i_0_26),
    .io_matrix_i_0_27(Reduction_2_io_matrix_i_0_27),
    .io_matrix_i_0_28(Reduction_2_io_matrix_i_0_28),
    .io_matrix_i_0_29(Reduction_2_io_matrix_i_0_29),
    .io_matrix_i_0_30(Reduction_2_io_matrix_i_0_30),
    .io_matrix_i_0_31(Reduction_2_io_matrix_i_0_31),
    .io_matrix_i_1_1(Reduction_2_io_matrix_i_1_1),
    .io_matrix_i_1_3(Reduction_2_io_matrix_i_1_3),
    .io_matrix_i_1_4(Reduction_2_io_matrix_i_1_4),
    .io_matrix_i_1_5(Reduction_2_io_matrix_i_1_5),
    .io_matrix_i_1_6(Reduction_2_io_matrix_i_1_6),
    .io_matrix_i_1_7(Reduction_2_io_matrix_i_1_7),
    .io_matrix_i_1_8(Reduction_2_io_matrix_i_1_8),
    .io_matrix_i_1_9(Reduction_2_io_matrix_i_1_9),
    .io_matrix_i_1_10(Reduction_2_io_matrix_i_1_10),
    .io_matrix_i_1_11(Reduction_2_io_matrix_i_1_11),
    .io_matrix_i_1_12(Reduction_2_io_matrix_i_1_12),
    .io_matrix_i_1_13(Reduction_2_io_matrix_i_1_13),
    .io_matrix_i_1_14(Reduction_2_io_matrix_i_1_14),
    .io_matrix_i_1_15(Reduction_2_io_matrix_i_1_15),
    .io_matrix_i_1_16(Reduction_2_io_matrix_i_1_16),
    .io_matrix_i_1_17(Reduction_2_io_matrix_i_1_17),
    .io_matrix_i_1_18(Reduction_2_io_matrix_i_1_18),
    .io_matrix_i_1_19(Reduction_2_io_matrix_i_1_19),
    .io_matrix_i_1_20(Reduction_2_io_matrix_i_1_20),
    .io_matrix_i_1_21(Reduction_2_io_matrix_i_1_21),
    .io_matrix_i_1_22(Reduction_2_io_matrix_i_1_22),
    .io_matrix_i_1_23(Reduction_2_io_matrix_i_1_23),
    .io_matrix_i_1_24(Reduction_2_io_matrix_i_1_24),
    .io_matrix_i_1_25(Reduction_2_io_matrix_i_1_25),
    .io_matrix_i_1_26(Reduction_2_io_matrix_i_1_26),
    .io_matrix_i_1_27(Reduction_2_io_matrix_i_1_27),
    .io_matrix_i_1_28(Reduction_2_io_matrix_i_1_28),
    .io_matrix_i_1_29(Reduction_2_io_matrix_i_1_29),
    .io_matrix_i_1_30(Reduction_2_io_matrix_i_1_30),
    .io_matrix_i_2_3(Reduction_2_io_matrix_i_2_3),
    .io_matrix_i_2_6(Reduction_2_io_matrix_i_2_6),
    .io_matrix_i_2_7(Reduction_2_io_matrix_i_2_7),
    .io_matrix_i_2_8(Reduction_2_io_matrix_i_2_8),
    .io_matrix_i_2_9(Reduction_2_io_matrix_i_2_9),
    .io_matrix_i_2_10(Reduction_2_io_matrix_i_2_10),
    .io_matrix_i_2_11(Reduction_2_io_matrix_i_2_11),
    .io_matrix_i_2_12(Reduction_2_io_matrix_i_2_12),
    .io_matrix_i_2_13(Reduction_2_io_matrix_i_2_13),
    .io_matrix_i_2_14(Reduction_2_io_matrix_i_2_14),
    .io_matrix_i_2_15(Reduction_2_io_matrix_i_2_15),
    .io_matrix_i_2_16(Reduction_2_io_matrix_i_2_16),
    .io_matrix_i_2_17(Reduction_2_io_matrix_i_2_17),
    .io_matrix_i_2_18(Reduction_2_io_matrix_i_2_18),
    .io_matrix_i_2_19(Reduction_2_io_matrix_i_2_19),
    .io_matrix_i_2_20(Reduction_2_io_matrix_i_2_20),
    .io_matrix_i_2_21(Reduction_2_io_matrix_i_2_21),
    .io_matrix_i_2_22(Reduction_2_io_matrix_i_2_22),
    .io_matrix_i_2_23(Reduction_2_io_matrix_i_2_23),
    .io_matrix_i_2_24(Reduction_2_io_matrix_i_2_24),
    .io_matrix_i_2_25(Reduction_2_io_matrix_i_2_25),
    .io_matrix_i_2_26(Reduction_2_io_matrix_i_2_26),
    .io_matrix_i_2_29(Reduction_2_io_matrix_i_2_29),
    .io_matrix_i_3_6(Reduction_2_io_matrix_i_3_6),
    .io_matrix_i_3_9(Reduction_2_io_matrix_i_3_9),
    .io_matrix_i_3_10(Reduction_2_io_matrix_i_3_10),
    .io_matrix_i_3_11(Reduction_2_io_matrix_i_3_11),
    .io_matrix_i_3_12(Reduction_2_io_matrix_i_3_12),
    .io_matrix_i_3_13(Reduction_2_io_matrix_i_3_13),
    .io_matrix_i_3_14(Reduction_2_io_matrix_i_3_14),
    .io_matrix_i_3_15(Reduction_2_io_matrix_i_3_15),
    .io_matrix_i_3_16(Reduction_2_io_matrix_i_3_16),
    .io_matrix_i_3_17(Reduction_2_io_matrix_i_3_17),
    .io_matrix_i_3_18(Reduction_2_io_matrix_i_3_18),
    .io_matrix_i_3_19(Reduction_2_io_matrix_i_3_19),
    .io_matrix_i_3_20(Reduction_2_io_matrix_i_3_20),
    .io_matrix_i_3_21(Reduction_2_io_matrix_i_3_21),
    .io_matrix_i_3_22(Reduction_2_io_matrix_i_3_22),
    .io_matrix_i_3_23(Reduction_2_io_matrix_i_3_23),
    .io_matrix_i_3_24(Reduction_2_io_matrix_i_3_24),
    .io_matrix_i_4_9(Reduction_2_io_matrix_i_4_9),
    .io_matrix_i_4_12(Reduction_2_io_matrix_i_4_12),
    .io_matrix_i_4_13(Reduction_2_io_matrix_i_4_13),
    .io_matrix_i_4_14(Reduction_2_io_matrix_i_4_14),
    .io_matrix_i_4_15(Reduction_2_io_matrix_i_4_15),
    .io_matrix_i_4_16(Reduction_2_io_matrix_i_4_16),
    .io_matrix_i_4_17(Reduction_2_io_matrix_i_4_17),
    .io_matrix_i_4_18(Reduction_2_io_matrix_i_4_18),
    .io_matrix_i_4_19(Reduction_2_io_matrix_i_4_19),
    .io_matrix_i_4_20(Reduction_2_io_matrix_i_4_20),
    .io_matrix_i_4_23(Reduction_2_io_matrix_i_4_23),
    .io_matrix_i_5_12(Reduction_2_io_matrix_i_5_12),
    .io_matrix_i_5_15(Reduction_2_io_matrix_i_5_15),
    .io_matrix_i_5_16(Reduction_2_io_matrix_i_5_16),
    .io_matrix_i_5_17(Reduction_2_io_matrix_i_5_17),
    .io_matrix_i_5_18(Reduction_2_io_matrix_i_5_18),
    .io_matrix_i_5_19(Reduction_2_io_matrix_i_5_19)
  );
  Reduction_3 Reduction_3 ( // @[RA_Mul.scala 535:21:@4753.4]
    .io_matrix_o_0_0(Reduction_3_io_matrix_o_0_0),
    .io_matrix_o_0_1(Reduction_3_io_matrix_o_0_1),
    .io_matrix_o_0_2(Reduction_3_io_matrix_o_0_2),
    .io_matrix_o_0_3(Reduction_3_io_matrix_o_0_3),
    .io_matrix_o_0_4(Reduction_3_io_matrix_o_0_4),
    .io_matrix_o_0_5(Reduction_3_io_matrix_o_0_5),
    .io_matrix_o_0_6(Reduction_3_io_matrix_o_0_6),
    .io_matrix_o_0_7(Reduction_3_io_matrix_o_0_7),
    .io_matrix_o_0_8(Reduction_3_io_matrix_o_0_8),
    .io_matrix_o_0_9(Reduction_3_io_matrix_o_0_9),
    .io_matrix_o_0_10(Reduction_3_io_matrix_o_0_10),
    .io_matrix_o_0_11(Reduction_3_io_matrix_o_0_11),
    .io_matrix_o_0_12(Reduction_3_io_matrix_o_0_12),
    .io_matrix_o_0_13(Reduction_3_io_matrix_o_0_13),
    .io_matrix_o_0_14(Reduction_3_io_matrix_o_0_14),
    .io_matrix_o_0_15(Reduction_3_io_matrix_o_0_15),
    .io_matrix_o_0_16(Reduction_3_io_matrix_o_0_16),
    .io_matrix_o_0_17(Reduction_3_io_matrix_o_0_17),
    .io_matrix_o_0_18(Reduction_3_io_matrix_o_0_18),
    .io_matrix_o_0_19(Reduction_3_io_matrix_o_0_19),
    .io_matrix_o_0_20(Reduction_3_io_matrix_o_0_20),
    .io_matrix_o_0_21(Reduction_3_io_matrix_o_0_21),
    .io_matrix_o_0_22(Reduction_3_io_matrix_o_0_22),
    .io_matrix_o_0_23(Reduction_3_io_matrix_o_0_23),
    .io_matrix_o_0_24(Reduction_3_io_matrix_o_0_24),
    .io_matrix_o_0_25(Reduction_3_io_matrix_o_0_25),
    .io_matrix_o_0_26(Reduction_3_io_matrix_o_0_26),
    .io_matrix_o_0_27(Reduction_3_io_matrix_o_0_27),
    .io_matrix_o_0_28(Reduction_3_io_matrix_o_0_28),
    .io_matrix_o_0_29(Reduction_3_io_matrix_o_0_29),
    .io_matrix_o_0_30(Reduction_3_io_matrix_o_0_30),
    .io_matrix_o_0_31(Reduction_3_io_matrix_o_0_31),
    .io_matrix_o_1_3(Reduction_3_io_matrix_o_1_3),
    .io_matrix_o_1_5(Reduction_3_io_matrix_o_1_5),
    .io_matrix_o_1_6(Reduction_3_io_matrix_o_1_6),
    .io_matrix_o_1_7(Reduction_3_io_matrix_o_1_7),
    .io_matrix_o_1_8(Reduction_3_io_matrix_o_1_8),
    .io_matrix_o_1_9(Reduction_3_io_matrix_o_1_9),
    .io_matrix_o_1_10(Reduction_3_io_matrix_o_1_10),
    .io_matrix_o_1_11(Reduction_3_io_matrix_o_1_11),
    .io_matrix_o_1_12(Reduction_3_io_matrix_o_1_12),
    .io_matrix_o_1_13(Reduction_3_io_matrix_o_1_13),
    .io_matrix_o_1_14(Reduction_3_io_matrix_o_1_14),
    .io_matrix_o_1_15(Reduction_3_io_matrix_o_1_15),
    .io_matrix_o_1_16(Reduction_3_io_matrix_o_1_16),
    .io_matrix_o_1_17(Reduction_3_io_matrix_o_1_17),
    .io_matrix_o_1_18(Reduction_3_io_matrix_o_1_18),
    .io_matrix_o_1_19(Reduction_3_io_matrix_o_1_19),
    .io_matrix_o_1_20(Reduction_3_io_matrix_o_1_20),
    .io_matrix_o_1_21(Reduction_3_io_matrix_o_1_21),
    .io_matrix_o_1_22(Reduction_3_io_matrix_o_1_22),
    .io_matrix_o_1_23(Reduction_3_io_matrix_o_1_23),
    .io_matrix_o_1_24(Reduction_3_io_matrix_o_1_24),
    .io_matrix_o_1_25(Reduction_3_io_matrix_o_1_25),
    .io_matrix_o_1_26(Reduction_3_io_matrix_o_1_26),
    .io_matrix_o_1_28(Reduction_3_io_matrix_o_1_28),
    .io_matrix_o_1_31(Reduction_3_io_matrix_o_1_31),
    .io_matrix_o_2_5(Reduction_3_io_matrix_o_2_5),
    .io_matrix_o_2_13(Reduction_3_io_matrix_o_2_13),
    .io_matrix_o_2_14(Reduction_3_io_matrix_o_2_14),
    .io_matrix_o_2_15(Reduction_3_io_matrix_o_2_15),
    .io_matrix_o_2_16(Reduction_3_io_matrix_o_2_16),
    .io_matrix_o_2_17(Reduction_3_io_matrix_o_2_17),
    .io_matrix_o_2_18(Reduction_3_io_matrix_o_2_18),
    .io_matrix_o_2_19(Reduction_3_io_matrix_o_2_19),
    .io_matrix_o_2_20(Reduction_3_io_matrix_o_2_20),
    .io_matrix_o_2_21(Reduction_3_io_matrix_o_2_21),
    .io_matrix_o_2_23(Reduction_3_io_matrix_o_2_23),
    .io_matrix_o_2_25(Reduction_3_io_matrix_o_2_25),
    .io_matrix_o_2_28(Reduction_3_io_matrix_o_2_28),
    .io_matrix_i_0_0(Reduction_3_io_matrix_i_0_0),
    .io_matrix_i_0_1(Reduction_3_io_matrix_i_0_1),
    .io_matrix_i_0_2(Reduction_3_io_matrix_i_0_2),
    .io_matrix_i_0_3(Reduction_3_io_matrix_i_0_3),
    .io_matrix_i_0_4(Reduction_3_io_matrix_i_0_4),
    .io_matrix_i_0_5(Reduction_3_io_matrix_i_0_5),
    .io_matrix_i_0_6(Reduction_3_io_matrix_i_0_6),
    .io_matrix_i_0_7(Reduction_3_io_matrix_i_0_7),
    .io_matrix_i_0_8(Reduction_3_io_matrix_i_0_8),
    .io_matrix_i_0_9(Reduction_3_io_matrix_i_0_9),
    .io_matrix_i_0_10(Reduction_3_io_matrix_i_0_10),
    .io_matrix_i_0_11(Reduction_3_io_matrix_i_0_11),
    .io_matrix_i_0_12(Reduction_3_io_matrix_i_0_12),
    .io_matrix_i_0_13(Reduction_3_io_matrix_i_0_13),
    .io_matrix_i_0_14(Reduction_3_io_matrix_i_0_14),
    .io_matrix_i_0_15(Reduction_3_io_matrix_i_0_15),
    .io_matrix_i_0_16(Reduction_3_io_matrix_i_0_16),
    .io_matrix_i_0_17(Reduction_3_io_matrix_i_0_17),
    .io_matrix_i_0_18(Reduction_3_io_matrix_i_0_18),
    .io_matrix_i_0_19(Reduction_3_io_matrix_i_0_19),
    .io_matrix_i_0_20(Reduction_3_io_matrix_i_0_20),
    .io_matrix_i_0_21(Reduction_3_io_matrix_i_0_21),
    .io_matrix_i_0_22(Reduction_3_io_matrix_i_0_22),
    .io_matrix_i_0_23(Reduction_3_io_matrix_i_0_23),
    .io_matrix_i_0_24(Reduction_3_io_matrix_i_0_24),
    .io_matrix_i_0_25(Reduction_3_io_matrix_i_0_25),
    .io_matrix_i_0_26(Reduction_3_io_matrix_i_0_26),
    .io_matrix_i_0_27(Reduction_3_io_matrix_i_0_27),
    .io_matrix_i_0_28(Reduction_3_io_matrix_i_0_28),
    .io_matrix_i_0_29(Reduction_3_io_matrix_i_0_29),
    .io_matrix_i_0_30(Reduction_3_io_matrix_i_0_30),
    .io_matrix_i_0_31(Reduction_3_io_matrix_i_0_31),
    .io_matrix_i_1_2(Reduction_3_io_matrix_i_1_2),
    .io_matrix_i_1_4(Reduction_3_io_matrix_i_1_4),
    .io_matrix_i_1_5(Reduction_3_io_matrix_i_1_5),
    .io_matrix_i_1_6(Reduction_3_io_matrix_i_1_6),
    .io_matrix_i_1_7(Reduction_3_io_matrix_i_1_7),
    .io_matrix_i_1_8(Reduction_3_io_matrix_i_1_8),
    .io_matrix_i_1_9(Reduction_3_io_matrix_i_1_9),
    .io_matrix_i_1_10(Reduction_3_io_matrix_i_1_10),
    .io_matrix_i_1_11(Reduction_3_io_matrix_i_1_11),
    .io_matrix_i_1_12(Reduction_3_io_matrix_i_1_12),
    .io_matrix_i_1_13(Reduction_3_io_matrix_i_1_13),
    .io_matrix_i_1_14(Reduction_3_io_matrix_i_1_14),
    .io_matrix_i_1_15(Reduction_3_io_matrix_i_1_15),
    .io_matrix_i_1_16(Reduction_3_io_matrix_i_1_16),
    .io_matrix_i_1_17(Reduction_3_io_matrix_i_1_17),
    .io_matrix_i_1_18(Reduction_3_io_matrix_i_1_18),
    .io_matrix_i_1_19(Reduction_3_io_matrix_i_1_19),
    .io_matrix_i_1_20(Reduction_3_io_matrix_i_1_20),
    .io_matrix_i_1_21(Reduction_3_io_matrix_i_1_21),
    .io_matrix_i_1_22(Reduction_3_io_matrix_i_1_22),
    .io_matrix_i_1_23(Reduction_3_io_matrix_i_1_23),
    .io_matrix_i_1_24(Reduction_3_io_matrix_i_1_24),
    .io_matrix_i_1_25(Reduction_3_io_matrix_i_1_25),
    .io_matrix_i_1_26(Reduction_3_io_matrix_i_1_26),
    .io_matrix_i_1_27(Reduction_3_io_matrix_i_1_27),
    .io_matrix_i_1_28(Reduction_3_io_matrix_i_1_28),
    .io_matrix_i_1_30(Reduction_3_io_matrix_i_1_30),
    .io_matrix_i_2_4(Reduction_3_io_matrix_i_2_4),
    .io_matrix_i_2_9(Reduction_3_io_matrix_i_2_9),
    .io_matrix_i_2_10(Reduction_3_io_matrix_i_2_10),
    .io_matrix_i_2_11(Reduction_3_io_matrix_i_2_11),
    .io_matrix_i_2_12(Reduction_3_io_matrix_i_2_12),
    .io_matrix_i_2_13(Reduction_3_io_matrix_i_2_13),
    .io_matrix_i_2_14(Reduction_3_io_matrix_i_2_14),
    .io_matrix_i_2_15(Reduction_3_io_matrix_i_2_15),
    .io_matrix_i_2_16(Reduction_3_io_matrix_i_2_16),
    .io_matrix_i_2_17(Reduction_3_io_matrix_i_2_17),
    .io_matrix_i_2_18(Reduction_3_io_matrix_i_2_18),
    .io_matrix_i_2_19(Reduction_3_io_matrix_i_2_19),
    .io_matrix_i_2_20(Reduction_3_io_matrix_i_2_20),
    .io_matrix_i_2_21(Reduction_3_io_matrix_i_2_21),
    .io_matrix_i_2_22(Reduction_3_io_matrix_i_2_22),
    .io_matrix_i_2_23(Reduction_3_io_matrix_i_2_23),
    .io_matrix_i_2_24(Reduction_3_io_matrix_i_2_24),
    .io_matrix_i_2_27(Reduction_3_io_matrix_i_2_27),
    .io_matrix_i_2_30(Reduction_3_io_matrix_i_2_30),
    .io_matrix_i_3_9(Reduction_3_io_matrix_i_3_9),
    .io_matrix_i_3_13(Reduction_3_io_matrix_i_3_13),
    .io_matrix_i_3_14(Reduction_3_io_matrix_i_3_14),
    .io_matrix_i_3_15(Reduction_3_io_matrix_i_3_15),
    .io_matrix_i_3_16(Reduction_3_io_matrix_i_3_16),
    .io_matrix_i_3_17(Reduction_3_io_matrix_i_3_17),
    .io_matrix_i_3_18(Reduction_3_io_matrix_i_3_18),
    .io_matrix_i_3_19(Reduction_3_io_matrix_i_3_19),
    .io_matrix_i_3_20(Reduction_3_io_matrix_i_3_20),
    .io_matrix_i_3_21(Reduction_3_io_matrix_i_3_21),
    .io_matrix_i_3_23(Reduction_3_io_matrix_i_3_23)
  );
  Reduction_4 Reduction_4 ( // @[RA_Mul.scala 598:21:@4980.4]
    .io_matrix_o_0_0(Reduction_4_io_matrix_o_0_0),
    .io_matrix_o_0_1(Reduction_4_io_matrix_o_0_1),
    .io_matrix_o_0_2(Reduction_4_io_matrix_o_0_2),
    .io_matrix_o_0_3(Reduction_4_io_matrix_o_0_3),
    .io_matrix_o_0_4(Reduction_4_io_matrix_o_0_4),
    .io_matrix_o_0_5(Reduction_4_io_matrix_o_0_5),
    .io_matrix_o_0_6(Reduction_4_io_matrix_o_0_6),
    .io_matrix_o_0_7(Reduction_4_io_matrix_o_0_7),
    .io_matrix_o_0_8(Reduction_4_io_matrix_o_0_8),
    .io_matrix_o_0_9(Reduction_4_io_matrix_o_0_9),
    .io_matrix_o_0_10(Reduction_4_io_matrix_o_0_10),
    .io_matrix_o_0_11(Reduction_4_io_matrix_o_0_11),
    .io_matrix_o_0_12(Reduction_4_io_matrix_o_0_12),
    .io_matrix_o_0_13(Reduction_4_io_matrix_o_0_13),
    .io_matrix_o_0_14(Reduction_4_io_matrix_o_0_14),
    .io_matrix_o_0_15(Reduction_4_io_matrix_o_0_15),
    .io_matrix_o_0_16(Reduction_4_io_matrix_o_0_16),
    .io_matrix_o_0_17(Reduction_4_io_matrix_o_0_17),
    .io_matrix_o_0_18(Reduction_4_io_matrix_o_0_18),
    .io_matrix_o_0_19(Reduction_4_io_matrix_o_0_19),
    .io_matrix_o_0_20(Reduction_4_io_matrix_o_0_20),
    .io_matrix_o_0_21(Reduction_4_io_matrix_o_0_21),
    .io_matrix_o_0_22(Reduction_4_io_matrix_o_0_22),
    .io_matrix_o_0_23(Reduction_4_io_matrix_o_0_23),
    .io_matrix_o_0_24(Reduction_4_io_matrix_o_0_24),
    .io_matrix_o_0_25(Reduction_4_io_matrix_o_0_25),
    .io_matrix_o_0_26(Reduction_4_io_matrix_o_0_26),
    .io_matrix_o_0_27(Reduction_4_io_matrix_o_0_27),
    .io_matrix_o_0_28(Reduction_4_io_matrix_o_0_28),
    .io_matrix_o_0_29(Reduction_4_io_matrix_o_0_29),
    .io_matrix_o_0_30(Reduction_4_io_matrix_o_0_30),
    .io_matrix_o_0_31(Reduction_4_io_matrix_o_0_31),
    .io_matrix_o_1_4(Reduction_4_io_matrix_o_1_4),
    .io_matrix_o_1_6(Reduction_4_io_matrix_o_1_6),
    .io_matrix_o_1_7(Reduction_4_io_matrix_o_1_7),
    .io_matrix_o_1_8(Reduction_4_io_matrix_o_1_8),
    .io_matrix_o_1_9(Reduction_4_io_matrix_o_1_9),
    .io_matrix_o_1_10(Reduction_4_io_matrix_o_1_10),
    .io_matrix_o_1_11(Reduction_4_io_matrix_o_1_11),
    .io_matrix_o_1_12(Reduction_4_io_matrix_o_1_12),
    .io_matrix_o_1_13(Reduction_4_io_matrix_o_1_13),
    .io_matrix_o_1_14(Reduction_4_io_matrix_o_1_14),
    .io_matrix_o_1_15(Reduction_4_io_matrix_o_1_15),
    .io_matrix_o_1_16(Reduction_4_io_matrix_o_1_16),
    .io_matrix_o_1_17(Reduction_4_io_matrix_o_1_17),
    .io_matrix_o_1_18(Reduction_4_io_matrix_o_1_18),
    .io_matrix_o_1_19(Reduction_4_io_matrix_o_1_19),
    .io_matrix_o_1_20(Reduction_4_io_matrix_o_1_20),
    .io_matrix_o_1_21(Reduction_4_io_matrix_o_1_21),
    .io_matrix_o_1_22(Reduction_4_io_matrix_o_1_22),
    .io_matrix_o_1_23(Reduction_4_io_matrix_o_1_23),
    .io_matrix_o_1_24(Reduction_4_io_matrix_o_1_24),
    .io_matrix_o_1_25(Reduction_4_io_matrix_o_1_25),
    .io_matrix_o_1_26(Reduction_4_io_matrix_o_1_26),
    .io_matrix_o_1_27(Reduction_4_io_matrix_o_1_27),
    .io_matrix_o_1_29(Reduction_4_io_matrix_o_1_29),
    .io_matrix_o_1_31(Reduction_4_io_matrix_o_1_31),
    .io_matrix_i_0_0(Reduction_4_io_matrix_i_0_0),
    .io_matrix_i_0_1(Reduction_4_io_matrix_i_0_1),
    .io_matrix_i_0_2(Reduction_4_io_matrix_i_0_2),
    .io_matrix_i_0_3(Reduction_4_io_matrix_i_0_3),
    .io_matrix_i_0_4(Reduction_4_io_matrix_i_0_4),
    .io_matrix_i_0_5(Reduction_4_io_matrix_i_0_5),
    .io_matrix_i_0_6(Reduction_4_io_matrix_i_0_6),
    .io_matrix_i_0_7(Reduction_4_io_matrix_i_0_7),
    .io_matrix_i_0_8(Reduction_4_io_matrix_i_0_8),
    .io_matrix_i_0_9(Reduction_4_io_matrix_i_0_9),
    .io_matrix_i_0_10(Reduction_4_io_matrix_i_0_10),
    .io_matrix_i_0_11(Reduction_4_io_matrix_i_0_11),
    .io_matrix_i_0_12(Reduction_4_io_matrix_i_0_12),
    .io_matrix_i_0_13(Reduction_4_io_matrix_i_0_13),
    .io_matrix_i_0_14(Reduction_4_io_matrix_i_0_14),
    .io_matrix_i_0_15(Reduction_4_io_matrix_i_0_15),
    .io_matrix_i_0_16(Reduction_4_io_matrix_i_0_16),
    .io_matrix_i_0_17(Reduction_4_io_matrix_i_0_17),
    .io_matrix_i_0_18(Reduction_4_io_matrix_i_0_18),
    .io_matrix_i_0_19(Reduction_4_io_matrix_i_0_19),
    .io_matrix_i_0_20(Reduction_4_io_matrix_i_0_20),
    .io_matrix_i_0_21(Reduction_4_io_matrix_i_0_21),
    .io_matrix_i_0_22(Reduction_4_io_matrix_i_0_22),
    .io_matrix_i_0_23(Reduction_4_io_matrix_i_0_23),
    .io_matrix_i_0_24(Reduction_4_io_matrix_i_0_24),
    .io_matrix_i_0_25(Reduction_4_io_matrix_i_0_25),
    .io_matrix_i_0_26(Reduction_4_io_matrix_i_0_26),
    .io_matrix_i_0_27(Reduction_4_io_matrix_i_0_27),
    .io_matrix_i_0_28(Reduction_4_io_matrix_i_0_28),
    .io_matrix_i_0_29(Reduction_4_io_matrix_i_0_29),
    .io_matrix_i_0_30(Reduction_4_io_matrix_i_0_30),
    .io_matrix_i_0_31(Reduction_4_io_matrix_i_0_31),
    .io_matrix_i_1_3(Reduction_4_io_matrix_i_1_3),
    .io_matrix_i_1_5(Reduction_4_io_matrix_i_1_5),
    .io_matrix_i_1_6(Reduction_4_io_matrix_i_1_6),
    .io_matrix_i_1_7(Reduction_4_io_matrix_i_1_7),
    .io_matrix_i_1_8(Reduction_4_io_matrix_i_1_8),
    .io_matrix_i_1_9(Reduction_4_io_matrix_i_1_9),
    .io_matrix_i_1_10(Reduction_4_io_matrix_i_1_10),
    .io_matrix_i_1_11(Reduction_4_io_matrix_i_1_11),
    .io_matrix_i_1_12(Reduction_4_io_matrix_i_1_12),
    .io_matrix_i_1_13(Reduction_4_io_matrix_i_1_13),
    .io_matrix_i_1_14(Reduction_4_io_matrix_i_1_14),
    .io_matrix_i_1_15(Reduction_4_io_matrix_i_1_15),
    .io_matrix_i_1_16(Reduction_4_io_matrix_i_1_16),
    .io_matrix_i_1_17(Reduction_4_io_matrix_i_1_17),
    .io_matrix_i_1_18(Reduction_4_io_matrix_i_1_18),
    .io_matrix_i_1_19(Reduction_4_io_matrix_i_1_19),
    .io_matrix_i_1_20(Reduction_4_io_matrix_i_1_20),
    .io_matrix_i_1_21(Reduction_4_io_matrix_i_1_21),
    .io_matrix_i_1_22(Reduction_4_io_matrix_i_1_22),
    .io_matrix_i_1_23(Reduction_4_io_matrix_i_1_23),
    .io_matrix_i_1_24(Reduction_4_io_matrix_i_1_24),
    .io_matrix_i_1_25(Reduction_4_io_matrix_i_1_25),
    .io_matrix_i_1_26(Reduction_4_io_matrix_i_1_26),
    .io_matrix_i_1_28(Reduction_4_io_matrix_i_1_28),
    .io_matrix_i_1_31(Reduction_4_io_matrix_i_1_31),
    .io_matrix_i_2_5(Reduction_4_io_matrix_i_2_5),
    .io_matrix_i_2_13(Reduction_4_io_matrix_i_2_13),
    .io_matrix_i_2_14(Reduction_4_io_matrix_i_2_14),
    .io_matrix_i_2_15(Reduction_4_io_matrix_i_2_15),
    .io_matrix_i_2_16(Reduction_4_io_matrix_i_2_16),
    .io_matrix_i_2_17(Reduction_4_io_matrix_i_2_17),
    .io_matrix_i_2_18(Reduction_4_io_matrix_i_2_18),
    .io_matrix_i_2_19(Reduction_4_io_matrix_i_2_19),
    .io_matrix_i_2_20(Reduction_4_io_matrix_i_2_20),
    .io_matrix_i_2_21(Reduction_4_io_matrix_i_2_21),
    .io_matrix_i_2_23(Reduction_4_io_matrix_i_2_23),
    .io_matrix_i_2_25(Reduction_4_io_matrix_i_2_25),
    .io_matrix_i_2_28(Reduction_4_io_matrix_i_2_28)
  );
  PPLRegs2 PPLRegs2 ( // @[RA_Mul.scala 711:21:@5143.4]
    .clock(PPLRegs2_clock),
    .reset(PPLRegs2_reset),
    .io_matrix_o_0_0(PPLRegs2_io_matrix_o_0_0),
    .io_matrix_o_0_1(PPLRegs2_io_matrix_o_0_1),
    .io_matrix_o_0_2(PPLRegs2_io_matrix_o_0_2),
    .io_matrix_o_0_3(PPLRegs2_io_matrix_o_0_3),
    .io_matrix_o_0_4(PPLRegs2_io_matrix_o_0_4),
    .io_matrix_o_0_5(PPLRegs2_io_matrix_o_0_5),
    .io_matrix_o_0_6(PPLRegs2_io_matrix_o_0_6),
    .io_matrix_o_0_7(PPLRegs2_io_matrix_o_0_7),
    .io_matrix_o_0_8(PPLRegs2_io_matrix_o_0_8),
    .io_matrix_o_0_9(PPLRegs2_io_matrix_o_0_9),
    .io_matrix_o_0_10(PPLRegs2_io_matrix_o_0_10),
    .io_matrix_o_0_11(PPLRegs2_io_matrix_o_0_11),
    .io_matrix_o_0_12(PPLRegs2_io_matrix_o_0_12),
    .io_matrix_o_0_13(PPLRegs2_io_matrix_o_0_13),
    .io_matrix_o_0_14(PPLRegs2_io_matrix_o_0_14),
    .io_matrix_o_0_15(PPLRegs2_io_matrix_o_0_15),
    .io_matrix_o_0_16(PPLRegs2_io_matrix_o_0_16),
    .io_matrix_o_0_17(PPLRegs2_io_matrix_o_0_17),
    .io_matrix_o_0_18(PPLRegs2_io_matrix_o_0_18),
    .io_matrix_o_0_19(PPLRegs2_io_matrix_o_0_19),
    .io_matrix_o_0_20(PPLRegs2_io_matrix_o_0_20),
    .io_matrix_o_0_21(PPLRegs2_io_matrix_o_0_21),
    .io_matrix_o_0_22(PPLRegs2_io_matrix_o_0_22),
    .io_matrix_o_0_23(PPLRegs2_io_matrix_o_0_23),
    .io_matrix_o_0_24(PPLRegs2_io_matrix_o_0_24),
    .io_matrix_o_0_25(PPLRegs2_io_matrix_o_0_25),
    .io_matrix_o_0_26(PPLRegs2_io_matrix_o_0_26),
    .io_matrix_o_0_27(PPLRegs2_io_matrix_o_0_27),
    .io_matrix_o_0_28(PPLRegs2_io_matrix_o_0_28),
    .io_matrix_o_0_29(PPLRegs2_io_matrix_o_0_29),
    .io_matrix_o_0_30(PPLRegs2_io_matrix_o_0_30),
    .io_matrix_o_0_31(PPLRegs2_io_matrix_o_0_31),
    .io_matrix_o_1_0(PPLRegs2_io_matrix_o_1_0),
    .io_matrix_o_1_1(PPLRegs2_io_matrix_o_1_1),
    .io_matrix_o_1_2(PPLRegs2_io_matrix_o_1_2),
    .io_matrix_o_1_3(PPLRegs2_io_matrix_o_1_3),
    .io_matrix_o_1_4(PPLRegs2_io_matrix_o_1_4),
    .io_matrix_o_1_5(PPLRegs2_io_matrix_o_1_5),
    .io_matrix_o_1_6(PPLRegs2_io_matrix_o_1_6),
    .io_matrix_o_1_7(PPLRegs2_io_matrix_o_1_7),
    .io_matrix_o_1_8(PPLRegs2_io_matrix_o_1_8),
    .io_matrix_o_1_9(PPLRegs2_io_matrix_o_1_9),
    .io_matrix_o_1_10(PPLRegs2_io_matrix_o_1_10),
    .io_matrix_o_1_11(PPLRegs2_io_matrix_o_1_11),
    .io_matrix_o_1_12(PPLRegs2_io_matrix_o_1_12),
    .io_matrix_o_1_13(PPLRegs2_io_matrix_o_1_13),
    .io_matrix_o_1_14(PPLRegs2_io_matrix_o_1_14),
    .io_matrix_o_1_15(PPLRegs2_io_matrix_o_1_15),
    .io_matrix_o_1_16(PPLRegs2_io_matrix_o_1_16),
    .io_matrix_o_1_17(PPLRegs2_io_matrix_o_1_17),
    .io_matrix_o_1_18(PPLRegs2_io_matrix_o_1_18),
    .io_matrix_o_1_19(PPLRegs2_io_matrix_o_1_19),
    .io_matrix_o_1_20(PPLRegs2_io_matrix_o_1_20),
    .io_matrix_o_1_21(PPLRegs2_io_matrix_o_1_21),
    .io_matrix_o_1_22(PPLRegs2_io_matrix_o_1_22),
    .io_matrix_o_1_23(PPLRegs2_io_matrix_o_1_23),
    .io_matrix_o_1_24(PPLRegs2_io_matrix_o_1_24),
    .io_matrix_o_1_25(PPLRegs2_io_matrix_o_1_25),
    .io_matrix_o_1_26(PPLRegs2_io_matrix_o_1_26),
    .io_matrix_o_1_27(PPLRegs2_io_matrix_o_1_27),
    .io_matrix_o_1_28(PPLRegs2_io_matrix_o_1_28),
    .io_matrix_o_1_29(PPLRegs2_io_matrix_o_1_29),
    .io_matrix_o_1_30(PPLRegs2_io_matrix_o_1_30),
    .io_matrix_o_1_31(PPLRegs2_io_matrix_o_1_31),
    .io_matrix_i_0_0(PPLRegs2_io_matrix_i_0_0),
    .io_matrix_i_0_1(PPLRegs2_io_matrix_i_0_1),
    .io_matrix_i_0_2(PPLRegs2_io_matrix_i_0_2),
    .io_matrix_i_0_3(PPLRegs2_io_matrix_i_0_3),
    .io_matrix_i_0_4(PPLRegs2_io_matrix_i_0_4),
    .io_matrix_i_0_5(PPLRegs2_io_matrix_i_0_5),
    .io_matrix_i_0_6(PPLRegs2_io_matrix_i_0_6),
    .io_matrix_i_0_7(PPLRegs2_io_matrix_i_0_7),
    .io_matrix_i_0_8(PPLRegs2_io_matrix_i_0_8),
    .io_matrix_i_0_9(PPLRegs2_io_matrix_i_0_9),
    .io_matrix_i_0_10(PPLRegs2_io_matrix_i_0_10),
    .io_matrix_i_0_11(PPLRegs2_io_matrix_i_0_11),
    .io_matrix_i_0_12(PPLRegs2_io_matrix_i_0_12),
    .io_matrix_i_0_13(PPLRegs2_io_matrix_i_0_13),
    .io_matrix_i_0_14(PPLRegs2_io_matrix_i_0_14),
    .io_matrix_i_0_15(PPLRegs2_io_matrix_i_0_15),
    .io_matrix_i_0_16(PPLRegs2_io_matrix_i_0_16),
    .io_matrix_i_0_17(PPLRegs2_io_matrix_i_0_17),
    .io_matrix_i_0_18(PPLRegs2_io_matrix_i_0_18),
    .io_matrix_i_0_19(PPLRegs2_io_matrix_i_0_19),
    .io_matrix_i_0_20(PPLRegs2_io_matrix_i_0_20),
    .io_matrix_i_0_21(PPLRegs2_io_matrix_i_0_21),
    .io_matrix_i_0_22(PPLRegs2_io_matrix_i_0_22),
    .io_matrix_i_0_23(PPLRegs2_io_matrix_i_0_23),
    .io_matrix_i_0_24(PPLRegs2_io_matrix_i_0_24),
    .io_matrix_i_0_25(PPLRegs2_io_matrix_i_0_25),
    .io_matrix_i_0_26(PPLRegs2_io_matrix_i_0_26),
    .io_matrix_i_0_27(PPLRegs2_io_matrix_i_0_27),
    .io_matrix_i_0_28(PPLRegs2_io_matrix_i_0_28),
    .io_matrix_i_0_29(PPLRegs2_io_matrix_i_0_29),
    .io_matrix_i_0_30(PPLRegs2_io_matrix_i_0_30),
    .io_matrix_i_0_31(PPLRegs2_io_matrix_i_0_31),
    .io_matrix_i_1_4(PPLRegs2_io_matrix_i_1_4),
    .io_matrix_i_1_6(PPLRegs2_io_matrix_i_1_6),
    .io_matrix_i_1_7(PPLRegs2_io_matrix_i_1_7),
    .io_matrix_i_1_8(PPLRegs2_io_matrix_i_1_8),
    .io_matrix_i_1_9(PPLRegs2_io_matrix_i_1_9),
    .io_matrix_i_1_10(PPLRegs2_io_matrix_i_1_10),
    .io_matrix_i_1_11(PPLRegs2_io_matrix_i_1_11),
    .io_matrix_i_1_12(PPLRegs2_io_matrix_i_1_12),
    .io_matrix_i_1_13(PPLRegs2_io_matrix_i_1_13),
    .io_matrix_i_1_14(PPLRegs2_io_matrix_i_1_14),
    .io_matrix_i_1_15(PPLRegs2_io_matrix_i_1_15),
    .io_matrix_i_1_16(PPLRegs2_io_matrix_i_1_16),
    .io_matrix_i_1_17(PPLRegs2_io_matrix_i_1_17),
    .io_matrix_i_1_18(PPLRegs2_io_matrix_i_1_18),
    .io_matrix_i_1_19(PPLRegs2_io_matrix_i_1_19),
    .io_matrix_i_1_20(PPLRegs2_io_matrix_i_1_20),
    .io_matrix_i_1_21(PPLRegs2_io_matrix_i_1_21),
    .io_matrix_i_1_22(PPLRegs2_io_matrix_i_1_22),
    .io_matrix_i_1_23(PPLRegs2_io_matrix_i_1_23),
    .io_matrix_i_1_24(PPLRegs2_io_matrix_i_1_24),
    .io_matrix_i_1_25(PPLRegs2_io_matrix_i_1_25),
    .io_matrix_i_1_26(PPLRegs2_io_matrix_i_1_26),
    .io_matrix_i_1_27(PPLRegs2_io_matrix_i_1_27),
    .io_matrix_i_1_29(PPLRegs2_io_matrix_i_1_29),
    .io_matrix_i_1_31(PPLRegs2_io_matrix_i_1_31)
  );
  TailAdder TailAdder ( // @[RA_Mul.scala 617:21:@5336.4]
    .io_S(TailAdder_io_S),
    .io_B(TailAdder_io_B),
    .io_A(TailAdder_io_A)
  );
  PPLRegs3 PPLRegs3 ( // @[RA_Mul.scala 729:21:@5342.4]
    .clock(PPLRegs3_clock),
    .reset(PPLRegs3_reset),
    .io_S_o(PPLRegs3_io_S_o),
    .io_S_i(PPLRegs3_io_S_i)
  );
  assign matrix_o4_o_0_1 = PPLRegs2_io_matrix_o_0_1; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5147.4]
  assign matrix_o4_o_0_0 = PPLRegs2_io_matrix_o_0_0; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5146.4]
  assign _T_3079 = {matrix_o4_o_0_1,matrix_o4_o_0_0}; // @[RA_Mul.scala 769:28:@5274.4]
  assign matrix_o4_o_0_3 = PPLRegs2_io_matrix_o_0_3; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5149.4]
  assign matrix_o4_o_0_2 = PPLRegs2_io_matrix_o_0_2; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5148.4]
  assign _T_3080 = {matrix_o4_o_0_3,matrix_o4_o_0_2}; // @[RA_Mul.scala 769:28:@5275.4]
  assign _T_3081 = {_T_3080,_T_3079}; // @[RA_Mul.scala 769:28:@5276.4]
  assign matrix_o4_o_0_5 = PPLRegs2_io_matrix_o_0_5; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5151.4]
  assign matrix_o4_o_0_4 = PPLRegs2_io_matrix_o_0_4; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5150.4]
  assign _T_3082 = {matrix_o4_o_0_5,matrix_o4_o_0_4}; // @[RA_Mul.scala 769:28:@5277.4]
  assign matrix_o4_o_0_7 = PPLRegs2_io_matrix_o_0_7; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5153.4]
  assign matrix_o4_o_0_6 = PPLRegs2_io_matrix_o_0_6; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5152.4]
  assign _T_3083 = {matrix_o4_o_0_7,matrix_o4_o_0_6}; // @[RA_Mul.scala 769:28:@5278.4]
  assign _T_3084 = {_T_3083,_T_3082}; // @[RA_Mul.scala 769:28:@5279.4]
  assign _T_3085 = {_T_3084,_T_3081}; // @[RA_Mul.scala 769:28:@5280.4]
  assign matrix_o4_o_0_9 = PPLRegs2_io_matrix_o_0_9; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5155.4]
  assign matrix_o4_o_0_8 = PPLRegs2_io_matrix_o_0_8; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5154.4]
  assign _T_3086 = {matrix_o4_o_0_9,matrix_o4_o_0_8}; // @[RA_Mul.scala 769:28:@5281.4]
  assign matrix_o4_o_0_11 = PPLRegs2_io_matrix_o_0_11; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5157.4]
  assign matrix_o4_o_0_10 = PPLRegs2_io_matrix_o_0_10; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5156.4]
  assign _T_3087 = {matrix_o4_o_0_11,matrix_o4_o_0_10}; // @[RA_Mul.scala 769:28:@5282.4]
  assign _T_3088 = {_T_3087,_T_3086}; // @[RA_Mul.scala 769:28:@5283.4]
  assign matrix_o4_o_0_13 = PPLRegs2_io_matrix_o_0_13; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5159.4]
  assign matrix_o4_o_0_12 = PPLRegs2_io_matrix_o_0_12; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5158.4]
  assign _T_3089 = {matrix_o4_o_0_13,matrix_o4_o_0_12}; // @[RA_Mul.scala 769:28:@5284.4]
  assign matrix_o4_o_0_15 = PPLRegs2_io_matrix_o_0_15; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5161.4]
  assign matrix_o4_o_0_14 = PPLRegs2_io_matrix_o_0_14; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5160.4]
  assign _T_3090 = {matrix_o4_o_0_15,matrix_o4_o_0_14}; // @[RA_Mul.scala 769:28:@5285.4]
  assign _T_3091 = {_T_3090,_T_3089}; // @[RA_Mul.scala 769:28:@5286.4]
  assign _T_3092 = {_T_3091,_T_3088}; // @[RA_Mul.scala 769:28:@5287.4]
  assign _T_3093 = {_T_3092,_T_3085}; // @[RA_Mul.scala 769:28:@5288.4]
  assign matrix_o4_o_0_17 = PPLRegs2_io_matrix_o_0_17; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5163.4]
  assign matrix_o4_o_0_16 = PPLRegs2_io_matrix_o_0_16; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5162.4]
  assign _T_3094 = {matrix_o4_o_0_17,matrix_o4_o_0_16}; // @[RA_Mul.scala 769:28:@5289.4]
  assign matrix_o4_o_0_19 = PPLRegs2_io_matrix_o_0_19; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5165.4]
  assign matrix_o4_o_0_18 = PPLRegs2_io_matrix_o_0_18; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5164.4]
  assign _T_3095 = {matrix_o4_o_0_19,matrix_o4_o_0_18}; // @[RA_Mul.scala 769:28:@5290.4]
  assign _T_3096 = {_T_3095,_T_3094}; // @[RA_Mul.scala 769:28:@5291.4]
  assign matrix_o4_o_0_21 = PPLRegs2_io_matrix_o_0_21; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5167.4]
  assign matrix_o4_o_0_20 = PPLRegs2_io_matrix_o_0_20; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5166.4]
  assign _T_3097 = {matrix_o4_o_0_21,matrix_o4_o_0_20}; // @[RA_Mul.scala 769:28:@5292.4]
  assign matrix_o4_o_0_23 = PPLRegs2_io_matrix_o_0_23; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5169.4]
  assign matrix_o4_o_0_22 = PPLRegs2_io_matrix_o_0_22; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5168.4]
  assign _T_3098 = {matrix_o4_o_0_23,matrix_o4_o_0_22}; // @[RA_Mul.scala 769:28:@5293.4]
  assign _T_3099 = {_T_3098,_T_3097}; // @[RA_Mul.scala 769:28:@5294.4]
  assign _T_3100 = {_T_3099,_T_3096}; // @[RA_Mul.scala 769:28:@5295.4]
  assign matrix_o4_o_0_25 = PPLRegs2_io_matrix_o_0_25; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5171.4]
  assign matrix_o4_o_0_24 = PPLRegs2_io_matrix_o_0_24; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5170.4]
  assign _T_3101 = {matrix_o4_o_0_25,matrix_o4_o_0_24}; // @[RA_Mul.scala 769:28:@5296.4]
  assign matrix_o4_o_0_27 = PPLRegs2_io_matrix_o_0_27; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5173.4]
  assign matrix_o4_o_0_26 = PPLRegs2_io_matrix_o_0_26; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5172.4]
  assign _T_3102 = {matrix_o4_o_0_27,matrix_o4_o_0_26}; // @[RA_Mul.scala 769:28:@5297.4]
  assign _T_3103 = {_T_3102,_T_3101}; // @[RA_Mul.scala 769:28:@5298.4]
  assign matrix_o4_o_0_29 = PPLRegs2_io_matrix_o_0_29; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5175.4]
  assign matrix_o4_o_0_28 = PPLRegs2_io_matrix_o_0_28; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5174.4]
  assign _T_3104 = {matrix_o4_o_0_29,matrix_o4_o_0_28}; // @[RA_Mul.scala 769:28:@5299.4]
  assign matrix_o4_o_0_31 = PPLRegs2_io_matrix_o_0_31; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5177.4]
  assign matrix_o4_o_0_30 = PPLRegs2_io_matrix_o_0_30; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5176.4]
  assign _T_3105 = {matrix_o4_o_0_31,matrix_o4_o_0_30}; // @[RA_Mul.scala 769:28:@5300.4]
  assign _T_3106 = {_T_3105,_T_3104}; // @[RA_Mul.scala 769:28:@5301.4]
  assign _T_3107 = {_T_3106,_T_3103}; // @[RA_Mul.scala 769:28:@5302.4]
  assign _T_3108 = {_T_3107,_T_3100}; // @[RA_Mul.scala 769:28:@5303.4]
  assign matrix_o4_o_1_1 = PPLRegs2_io_matrix_o_1_1; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5179.4]
  assign matrix_o4_o_1_0 = PPLRegs2_io_matrix_o_1_0; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5178.4]
  assign _T_3110 = {matrix_o4_o_1_1,matrix_o4_o_1_0}; // @[RA_Mul.scala 769:51:@5305.4]
  assign matrix_o4_o_1_3 = PPLRegs2_io_matrix_o_1_3; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5181.4]
  assign matrix_o4_o_1_2 = PPLRegs2_io_matrix_o_1_2; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5180.4]
  assign _T_3111 = {matrix_o4_o_1_3,matrix_o4_o_1_2}; // @[RA_Mul.scala 769:51:@5306.4]
  assign _T_3112 = {_T_3111,_T_3110}; // @[RA_Mul.scala 769:51:@5307.4]
  assign matrix_o4_o_1_5 = PPLRegs2_io_matrix_o_1_5; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5183.4]
  assign matrix_o4_o_1_4 = PPLRegs2_io_matrix_o_1_4; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5182.4]
  assign _T_3113 = {matrix_o4_o_1_5,matrix_o4_o_1_4}; // @[RA_Mul.scala 769:51:@5308.4]
  assign matrix_o4_o_1_7 = PPLRegs2_io_matrix_o_1_7; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5185.4]
  assign matrix_o4_o_1_6 = PPLRegs2_io_matrix_o_1_6; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5184.4]
  assign _T_3114 = {matrix_o4_o_1_7,matrix_o4_o_1_6}; // @[RA_Mul.scala 769:51:@5309.4]
  assign _T_3115 = {_T_3114,_T_3113}; // @[RA_Mul.scala 769:51:@5310.4]
  assign _T_3116 = {_T_3115,_T_3112}; // @[RA_Mul.scala 769:51:@5311.4]
  assign matrix_o4_o_1_9 = PPLRegs2_io_matrix_o_1_9; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5187.4]
  assign matrix_o4_o_1_8 = PPLRegs2_io_matrix_o_1_8; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5186.4]
  assign _T_3117 = {matrix_o4_o_1_9,matrix_o4_o_1_8}; // @[RA_Mul.scala 769:51:@5312.4]
  assign matrix_o4_o_1_11 = PPLRegs2_io_matrix_o_1_11; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5189.4]
  assign matrix_o4_o_1_10 = PPLRegs2_io_matrix_o_1_10; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5188.4]
  assign _T_3118 = {matrix_o4_o_1_11,matrix_o4_o_1_10}; // @[RA_Mul.scala 769:51:@5313.4]
  assign _T_3119 = {_T_3118,_T_3117}; // @[RA_Mul.scala 769:51:@5314.4]
  assign matrix_o4_o_1_13 = PPLRegs2_io_matrix_o_1_13; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5191.4]
  assign matrix_o4_o_1_12 = PPLRegs2_io_matrix_o_1_12; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5190.4]
  assign _T_3120 = {matrix_o4_o_1_13,matrix_o4_o_1_12}; // @[RA_Mul.scala 769:51:@5315.4]
  assign matrix_o4_o_1_15 = PPLRegs2_io_matrix_o_1_15; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5193.4]
  assign matrix_o4_o_1_14 = PPLRegs2_io_matrix_o_1_14; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5192.4]
  assign _T_3121 = {matrix_o4_o_1_15,matrix_o4_o_1_14}; // @[RA_Mul.scala 769:51:@5316.4]
  assign _T_3122 = {_T_3121,_T_3120}; // @[RA_Mul.scala 769:51:@5317.4]
  assign _T_3123 = {_T_3122,_T_3119}; // @[RA_Mul.scala 769:51:@5318.4]
  assign _T_3124 = {_T_3123,_T_3116}; // @[RA_Mul.scala 769:51:@5319.4]
  assign matrix_o4_o_1_17 = PPLRegs2_io_matrix_o_1_17; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5195.4]
  assign matrix_o4_o_1_16 = PPLRegs2_io_matrix_o_1_16; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5194.4]
  assign _T_3125 = {matrix_o4_o_1_17,matrix_o4_o_1_16}; // @[RA_Mul.scala 769:51:@5320.4]
  assign matrix_o4_o_1_19 = PPLRegs2_io_matrix_o_1_19; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5197.4]
  assign matrix_o4_o_1_18 = PPLRegs2_io_matrix_o_1_18; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5196.4]
  assign _T_3126 = {matrix_o4_o_1_19,matrix_o4_o_1_18}; // @[RA_Mul.scala 769:51:@5321.4]
  assign _T_3127 = {_T_3126,_T_3125}; // @[RA_Mul.scala 769:51:@5322.4]
  assign matrix_o4_o_1_21 = PPLRegs2_io_matrix_o_1_21; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5199.4]
  assign matrix_o4_o_1_20 = PPLRegs2_io_matrix_o_1_20; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5198.4]
  assign _T_3128 = {matrix_o4_o_1_21,matrix_o4_o_1_20}; // @[RA_Mul.scala 769:51:@5323.4]
  assign matrix_o4_o_1_23 = PPLRegs2_io_matrix_o_1_23; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5201.4]
  assign matrix_o4_o_1_22 = PPLRegs2_io_matrix_o_1_22; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5200.4]
  assign _T_3129 = {matrix_o4_o_1_23,matrix_o4_o_1_22}; // @[RA_Mul.scala 769:51:@5324.4]
  assign _T_3130 = {_T_3129,_T_3128}; // @[RA_Mul.scala 769:51:@5325.4]
  assign _T_3131 = {_T_3130,_T_3127}; // @[RA_Mul.scala 769:51:@5326.4]
  assign matrix_o4_o_1_25 = PPLRegs2_io_matrix_o_1_25; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5203.4]
  assign matrix_o4_o_1_24 = PPLRegs2_io_matrix_o_1_24; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5202.4]
  assign _T_3132 = {matrix_o4_o_1_25,matrix_o4_o_1_24}; // @[RA_Mul.scala 769:51:@5327.4]
  assign matrix_o4_o_1_27 = PPLRegs2_io_matrix_o_1_27; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5205.4]
  assign matrix_o4_o_1_26 = PPLRegs2_io_matrix_o_1_26; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5204.4]
  assign _T_3133 = {matrix_o4_o_1_27,matrix_o4_o_1_26}; // @[RA_Mul.scala 769:51:@5328.4]
  assign _T_3134 = {_T_3133,_T_3132}; // @[RA_Mul.scala 769:51:@5329.4]
  assign matrix_o4_o_1_29 = PPLRegs2_io_matrix_o_1_29; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5207.4]
  assign matrix_o4_o_1_28 = PPLRegs2_io_matrix_o_1_28; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5206.4]
  assign _T_3135 = {matrix_o4_o_1_29,matrix_o4_o_1_28}; // @[RA_Mul.scala 769:51:@5330.4]
  assign matrix_o4_o_1_31 = PPLRegs2_io_matrix_o_1_31; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5209.4]
  assign matrix_o4_o_1_30 = PPLRegs2_io_matrix_o_1_30; // @[RA_Mul.scala 756:25:@4162.4 RA_Mul.scala 713:9:@5208.4]
  assign _T_3136 = {matrix_o4_o_1_31,matrix_o4_o_1_30}; // @[RA_Mul.scala 769:51:@5331.4]
  assign _T_3137 = {_T_3136,_T_3135}; // @[RA_Mul.scala 769:51:@5332.4]
  assign _T_3138 = {_T_3137,_T_3134}; // @[RA_Mul.scala 769:51:@5333.4]
  assign _T_3139 = {_T_3138,_T_3131}; // @[RA_Mul.scala 769:51:@5334.4]
  assign io_P = PPLRegs3_io_S_o; // @[RA_Mul.scala 731:9:@5346.4]
  assign BoothEncoder_radix4_io_B = io_B; // @[RA_Mul.scala 106:14:@4167.4]
  assign PPGen_io_eB_0 = BoothEncoder_radix4_io_eB_0; // @[RA_Mul.scala 161:15:@4180.4]
  assign PPGen_io_eB_1 = BoothEncoder_radix4_io_eB_1; // @[RA_Mul.scala 161:15:@4181.4]
  assign PPGen_io_eB_2 = BoothEncoder_radix4_io_eB_2; // @[RA_Mul.scala 161:15:@4182.4]
  assign PPGen_io_eB_3 = BoothEncoder_radix4_io_eB_3; // @[RA_Mul.scala 161:15:@4183.4]
  assign PPGen_io_eB_4 = BoothEncoder_radix4_io_eB_4; // @[RA_Mul.scala 161:15:@4184.4]
  assign PPGen_io_eB_5 = BoothEncoder_radix4_io_eB_5; // @[RA_Mul.scala 161:15:@4185.4]
  assign PPGen_io_eB_6 = BoothEncoder_radix4_io_eB_6; // @[RA_Mul.scala 161:15:@4186.4]
  assign PPGen_io_eB_7 = BoothEncoder_radix4_io_eB_7; // @[RA_Mul.scala 161:15:@4187.4]
  assign PPGen_io_A = io_A; // @[RA_Mul.scala 160:14:@4179.4]
  assign PPLRegs1_clock = clock; // @[:@4200.4]
  assign PPLRegs1_reset = reset; // @[:@4201.4]
  assign PPLRegs1_io_PP_i_0 = PPGen_io_PP_0; // @[RA_Mul.scala 680:17:@4202.4]
  assign PPLRegs1_io_PP_i_1 = PPGen_io_PP_1; // @[RA_Mul.scala 680:17:@4203.4]
  assign PPLRegs1_io_PP_i_2 = PPGen_io_PP_2; // @[RA_Mul.scala 680:17:@4204.4]
  assign PPLRegs1_io_PP_i_3 = PPGen_io_PP_3; // @[RA_Mul.scala 680:17:@4205.4]
  assign PPLRegs1_io_PP_i_4 = PPGen_io_PP_4; // @[RA_Mul.scala 680:17:@4206.4]
  assign PPLRegs1_io_PP_i_5 = PPGen_io_PP_5; // @[RA_Mul.scala 680:17:@4207.4]
  assign PPLRegs1_io_PP_i_6 = PPGen_io_PP_6; // @[RA_Mul.scala 680:17:@4208.4]
  assign PPLRegs1_io_PP_i_7 = PPGen_io_PP_7; // @[RA_Mul.scala 680:17:@4209.4]
  assign PPLRegs1_io_SC_i = PPGen_io_SC; // @[RA_Mul.scala 686:17:@4220.4]
  assign PPLRegs1_io_S_i = PPGen_io_S; // @[RA_Mul.scala 688:16:@4222.4]
  assign Reduction_1_io_PP_0 = PPLRegs1_io_PP_o_0; // @[RA_Mul.scala 321:15:@4227.4]
  assign Reduction_1_io_PP_1 = PPLRegs1_io_PP_o_1; // @[RA_Mul.scala 321:15:@4228.4]
  assign Reduction_1_io_PP_2 = PPLRegs1_io_PP_o_2; // @[RA_Mul.scala 321:15:@4229.4]
  assign Reduction_1_io_PP_3 = PPLRegs1_io_PP_o_3; // @[RA_Mul.scala 321:15:@4230.4]
  assign Reduction_1_io_PP_4 = PPLRegs1_io_PP_o_4; // @[RA_Mul.scala 321:15:@4231.4]
  assign Reduction_1_io_PP_5 = PPLRegs1_io_PP_o_5; // @[RA_Mul.scala 321:15:@4232.4]
  assign Reduction_1_io_PP_6 = PPLRegs1_io_PP_o_6; // @[RA_Mul.scala 321:15:@4233.4]
  assign Reduction_1_io_PP_7 = PPLRegs1_io_PP_o_7; // @[RA_Mul.scala 321:15:@4234.4]
  assign Reduction_1_io_SS = PPLRegs1_io_SS_o; // @[RA_Mul.scala 322:15:@4235.4]
  assign Reduction_1_io_SC = PPLRegs1_io_SC_o; // @[RA_Mul.scala 323:15:@4236.4]
  assign Reduction_1_io_S = PPLRegs1_io_S_o; // @[RA_Mul.scala 324:14:@4237.4]
  assign Reduction_2_io_matrix_i_0_0 = Reduction_1_io_matrix_0_0; // @[RA_Mul.scala 446:9:@4433.4]
  assign Reduction_2_io_matrix_i_0_1 = Reduction_1_io_matrix_0_1; // @[RA_Mul.scala 446:9:@4434.4]
  assign Reduction_2_io_matrix_i_0_2 = Reduction_1_io_matrix_0_2; // @[RA_Mul.scala 446:9:@4435.4]
  assign Reduction_2_io_matrix_i_0_3 = Reduction_1_io_matrix_0_3; // @[RA_Mul.scala 446:9:@4436.4]
  assign Reduction_2_io_matrix_i_0_4 = Reduction_1_io_matrix_0_4; // @[RA_Mul.scala 446:9:@4437.4]
  assign Reduction_2_io_matrix_i_0_5 = Reduction_1_io_matrix_0_5; // @[RA_Mul.scala 446:9:@4438.4]
  assign Reduction_2_io_matrix_i_0_6 = Reduction_1_io_matrix_0_6; // @[RA_Mul.scala 446:9:@4439.4]
  assign Reduction_2_io_matrix_i_0_7 = Reduction_1_io_matrix_0_7; // @[RA_Mul.scala 446:9:@4440.4]
  assign Reduction_2_io_matrix_i_0_8 = Reduction_1_io_matrix_0_8; // @[RA_Mul.scala 446:9:@4441.4]
  assign Reduction_2_io_matrix_i_0_9 = Reduction_1_io_matrix_0_9; // @[RA_Mul.scala 446:9:@4442.4]
  assign Reduction_2_io_matrix_i_0_10 = Reduction_1_io_matrix_0_10; // @[RA_Mul.scala 446:9:@4443.4]
  assign Reduction_2_io_matrix_i_0_11 = Reduction_1_io_matrix_0_11; // @[RA_Mul.scala 446:9:@4444.4]
  assign Reduction_2_io_matrix_i_0_12 = Reduction_1_io_matrix_0_12; // @[RA_Mul.scala 446:9:@4445.4]
  assign Reduction_2_io_matrix_i_0_13 = Reduction_1_io_matrix_0_13; // @[RA_Mul.scala 446:9:@4446.4]
  assign Reduction_2_io_matrix_i_0_14 = Reduction_1_io_matrix_0_14; // @[RA_Mul.scala 446:9:@4447.4]
  assign Reduction_2_io_matrix_i_0_15 = Reduction_1_io_matrix_0_15; // @[RA_Mul.scala 446:9:@4448.4]
  assign Reduction_2_io_matrix_i_0_16 = Reduction_1_io_matrix_0_16; // @[RA_Mul.scala 446:9:@4449.4]
  assign Reduction_2_io_matrix_i_0_17 = Reduction_1_io_matrix_0_17; // @[RA_Mul.scala 446:9:@4450.4]
  assign Reduction_2_io_matrix_i_0_18 = Reduction_1_io_matrix_0_18; // @[RA_Mul.scala 446:9:@4451.4]
  assign Reduction_2_io_matrix_i_0_19 = Reduction_1_io_matrix_0_19; // @[RA_Mul.scala 446:9:@4452.4]
  assign Reduction_2_io_matrix_i_0_20 = Reduction_1_io_matrix_0_20; // @[RA_Mul.scala 446:9:@4453.4]
  assign Reduction_2_io_matrix_i_0_21 = Reduction_1_io_matrix_0_21; // @[RA_Mul.scala 446:9:@4454.4]
  assign Reduction_2_io_matrix_i_0_22 = Reduction_1_io_matrix_0_22; // @[RA_Mul.scala 446:9:@4455.4]
  assign Reduction_2_io_matrix_i_0_23 = Reduction_1_io_matrix_0_23; // @[RA_Mul.scala 446:9:@4456.4]
  assign Reduction_2_io_matrix_i_0_24 = Reduction_1_io_matrix_0_24; // @[RA_Mul.scala 446:9:@4457.4]
  assign Reduction_2_io_matrix_i_0_25 = Reduction_1_io_matrix_0_25; // @[RA_Mul.scala 446:9:@4458.4]
  assign Reduction_2_io_matrix_i_0_26 = Reduction_1_io_matrix_0_26; // @[RA_Mul.scala 446:9:@4459.4]
  assign Reduction_2_io_matrix_i_0_27 = Reduction_1_io_matrix_0_27; // @[RA_Mul.scala 446:9:@4460.4]
  assign Reduction_2_io_matrix_i_0_28 = Reduction_1_io_matrix_0_28; // @[RA_Mul.scala 446:9:@4461.4]
  assign Reduction_2_io_matrix_i_0_29 = Reduction_1_io_matrix_0_29; // @[RA_Mul.scala 446:9:@4462.4]
  assign Reduction_2_io_matrix_i_0_30 = Reduction_1_io_matrix_0_30; // @[RA_Mul.scala 446:9:@4463.4]
  assign Reduction_2_io_matrix_i_0_31 = Reduction_1_io_matrix_0_31; // @[RA_Mul.scala 446:9:@4464.4]
  assign Reduction_2_io_matrix_i_1_1 = Reduction_1_io_matrix_1_1; // @[RA_Mul.scala 446:9:@4466.4]
  assign Reduction_2_io_matrix_i_1_3 = Reduction_1_io_matrix_1_3; // @[RA_Mul.scala 446:9:@4468.4]
  assign Reduction_2_io_matrix_i_1_4 = Reduction_1_io_matrix_1_4; // @[RA_Mul.scala 446:9:@4469.4]
  assign Reduction_2_io_matrix_i_1_5 = Reduction_1_io_matrix_1_5; // @[RA_Mul.scala 446:9:@4470.4]
  assign Reduction_2_io_matrix_i_1_6 = Reduction_1_io_matrix_1_6; // @[RA_Mul.scala 446:9:@4471.4]
  assign Reduction_2_io_matrix_i_1_7 = Reduction_1_io_matrix_1_7; // @[RA_Mul.scala 446:9:@4472.4]
  assign Reduction_2_io_matrix_i_1_8 = Reduction_1_io_matrix_1_8; // @[RA_Mul.scala 446:9:@4473.4]
  assign Reduction_2_io_matrix_i_1_9 = Reduction_1_io_matrix_1_9; // @[RA_Mul.scala 446:9:@4474.4]
  assign Reduction_2_io_matrix_i_1_10 = Reduction_1_io_matrix_1_10; // @[RA_Mul.scala 446:9:@4475.4]
  assign Reduction_2_io_matrix_i_1_11 = Reduction_1_io_matrix_1_11; // @[RA_Mul.scala 446:9:@4476.4]
  assign Reduction_2_io_matrix_i_1_12 = Reduction_1_io_matrix_1_12; // @[RA_Mul.scala 446:9:@4477.4]
  assign Reduction_2_io_matrix_i_1_13 = Reduction_1_io_matrix_1_13; // @[RA_Mul.scala 446:9:@4478.4]
  assign Reduction_2_io_matrix_i_1_14 = Reduction_1_io_matrix_1_14; // @[RA_Mul.scala 446:9:@4479.4]
  assign Reduction_2_io_matrix_i_1_15 = Reduction_1_io_matrix_1_15; // @[RA_Mul.scala 446:9:@4480.4]
  assign Reduction_2_io_matrix_i_1_16 = Reduction_1_io_matrix_1_16; // @[RA_Mul.scala 446:9:@4481.4]
  assign Reduction_2_io_matrix_i_1_17 = Reduction_1_io_matrix_1_17; // @[RA_Mul.scala 446:9:@4482.4]
  assign Reduction_2_io_matrix_i_1_18 = Reduction_1_io_matrix_1_18; // @[RA_Mul.scala 446:9:@4483.4]
  assign Reduction_2_io_matrix_i_1_19 = Reduction_1_io_matrix_1_19; // @[RA_Mul.scala 446:9:@4484.4]
  assign Reduction_2_io_matrix_i_1_20 = Reduction_1_io_matrix_1_20; // @[RA_Mul.scala 446:9:@4485.4]
  assign Reduction_2_io_matrix_i_1_21 = Reduction_1_io_matrix_1_21; // @[RA_Mul.scala 446:9:@4486.4]
  assign Reduction_2_io_matrix_i_1_22 = Reduction_1_io_matrix_1_22; // @[RA_Mul.scala 446:9:@4487.4]
  assign Reduction_2_io_matrix_i_1_23 = Reduction_1_io_matrix_1_23; // @[RA_Mul.scala 446:9:@4488.4]
  assign Reduction_2_io_matrix_i_1_24 = Reduction_1_io_matrix_1_24; // @[RA_Mul.scala 446:9:@4489.4]
  assign Reduction_2_io_matrix_i_1_25 = Reduction_1_io_matrix_1_25; // @[RA_Mul.scala 446:9:@4490.4]
  assign Reduction_2_io_matrix_i_1_26 = Reduction_1_io_matrix_1_26; // @[RA_Mul.scala 446:9:@4491.4]
  assign Reduction_2_io_matrix_i_1_27 = Reduction_1_io_matrix_1_27; // @[RA_Mul.scala 446:9:@4492.4]
  assign Reduction_2_io_matrix_i_1_28 = Reduction_1_io_matrix_1_28; // @[RA_Mul.scala 446:9:@4493.4]
  assign Reduction_2_io_matrix_i_1_29 = Reduction_1_io_matrix_1_29; // @[RA_Mul.scala 446:9:@4494.4]
  assign Reduction_2_io_matrix_i_1_30 = Reduction_1_io_matrix_1_30; // @[RA_Mul.scala 446:9:@4495.4]
  assign Reduction_2_io_matrix_i_2_3 = Reduction_1_io_matrix_2_3; // @[RA_Mul.scala 446:9:@4500.4]
  assign Reduction_2_io_matrix_i_2_6 = Reduction_1_io_matrix_2_6; // @[RA_Mul.scala 446:9:@4503.4]
  assign Reduction_2_io_matrix_i_2_7 = Reduction_1_io_matrix_2_7; // @[RA_Mul.scala 446:9:@4504.4]
  assign Reduction_2_io_matrix_i_2_8 = Reduction_1_io_matrix_2_8; // @[RA_Mul.scala 446:9:@4505.4]
  assign Reduction_2_io_matrix_i_2_9 = Reduction_1_io_matrix_2_9; // @[RA_Mul.scala 446:9:@4506.4]
  assign Reduction_2_io_matrix_i_2_10 = Reduction_1_io_matrix_2_10; // @[RA_Mul.scala 446:9:@4507.4]
  assign Reduction_2_io_matrix_i_2_11 = Reduction_1_io_matrix_2_11; // @[RA_Mul.scala 446:9:@4508.4]
  assign Reduction_2_io_matrix_i_2_12 = Reduction_1_io_matrix_2_12; // @[RA_Mul.scala 446:9:@4509.4]
  assign Reduction_2_io_matrix_i_2_13 = Reduction_1_io_matrix_2_13; // @[RA_Mul.scala 446:9:@4510.4]
  assign Reduction_2_io_matrix_i_2_14 = Reduction_1_io_matrix_2_14; // @[RA_Mul.scala 446:9:@4511.4]
  assign Reduction_2_io_matrix_i_2_15 = Reduction_1_io_matrix_2_15; // @[RA_Mul.scala 446:9:@4512.4]
  assign Reduction_2_io_matrix_i_2_16 = Reduction_1_io_matrix_2_16; // @[RA_Mul.scala 446:9:@4513.4]
  assign Reduction_2_io_matrix_i_2_17 = Reduction_1_io_matrix_2_17; // @[RA_Mul.scala 446:9:@4514.4]
  assign Reduction_2_io_matrix_i_2_18 = Reduction_1_io_matrix_2_18; // @[RA_Mul.scala 446:9:@4515.4]
  assign Reduction_2_io_matrix_i_2_19 = Reduction_1_io_matrix_2_19; // @[RA_Mul.scala 446:9:@4516.4]
  assign Reduction_2_io_matrix_i_2_20 = Reduction_1_io_matrix_2_20; // @[RA_Mul.scala 446:9:@4517.4]
  assign Reduction_2_io_matrix_i_2_21 = Reduction_1_io_matrix_2_21; // @[RA_Mul.scala 446:9:@4518.4]
  assign Reduction_2_io_matrix_i_2_22 = Reduction_1_io_matrix_2_22; // @[RA_Mul.scala 446:9:@4519.4]
  assign Reduction_2_io_matrix_i_2_23 = Reduction_1_io_matrix_2_23; // @[RA_Mul.scala 446:9:@4520.4]
  assign Reduction_2_io_matrix_i_2_24 = Reduction_1_io_matrix_2_24; // @[RA_Mul.scala 446:9:@4521.4]
  assign Reduction_2_io_matrix_i_2_25 = Reduction_1_io_matrix_2_25; // @[RA_Mul.scala 446:9:@4522.4]
  assign Reduction_2_io_matrix_i_2_26 = Reduction_1_io_matrix_2_26; // @[RA_Mul.scala 446:9:@4523.4]
  assign Reduction_2_io_matrix_i_2_29 = Reduction_1_io_matrix_2_29; // @[RA_Mul.scala 446:9:@4526.4]
  assign Reduction_2_io_matrix_i_3_6 = Reduction_1_io_matrix_3_6; // @[RA_Mul.scala 446:9:@4535.4]
  assign Reduction_2_io_matrix_i_3_9 = Reduction_1_io_matrix_3_9; // @[RA_Mul.scala 446:9:@4538.4]
  assign Reduction_2_io_matrix_i_3_10 = Reduction_1_io_matrix_3_10; // @[RA_Mul.scala 446:9:@4539.4]
  assign Reduction_2_io_matrix_i_3_11 = Reduction_1_io_matrix_3_11; // @[RA_Mul.scala 446:9:@4540.4]
  assign Reduction_2_io_matrix_i_3_12 = Reduction_1_io_matrix_3_12; // @[RA_Mul.scala 446:9:@4541.4]
  assign Reduction_2_io_matrix_i_3_13 = Reduction_1_io_matrix_3_13; // @[RA_Mul.scala 446:9:@4542.4]
  assign Reduction_2_io_matrix_i_3_14 = Reduction_1_io_matrix_3_14; // @[RA_Mul.scala 446:9:@4543.4]
  assign Reduction_2_io_matrix_i_3_15 = Reduction_1_io_matrix_3_15; // @[RA_Mul.scala 446:9:@4544.4]
  assign Reduction_2_io_matrix_i_3_16 = Reduction_1_io_matrix_3_16; // @[RA_Mul.scala 446:9:@4545.4]
  assign Reduction_2_io_matrix_i_3_17 = Reduction_1_io_matrix_3_17; // @[RA_Mul.scala 446:9:@4546.4]
  assign Reduction_2_io_matrix_i_3_18 = Reduction_1_io_matrix_3_18; // @[RA_Mul.scala 446:9:@4547.4]
  assign Reduction_2_io_matrix_i_3_19 = Reduction_1_io_matrix_3_19; // @[RA_Mul.scala 446:9:@4548.4]
  assign Reduction_2_io_matrix_i_3_20 = Reduction_1_io_matrix_3_20; // @[RA_Mul.scala 446:9:@4549.4]
  assign Reduction_2_io_matrix_i_3_21 = Reduction_1_io_matrix_3_21; // @[RA_Mul.scala 446:9:@4550.4]
  assign Reduction_2_io_matrix_i_3_22 = Reduction_1_io_matrix_3_22; // @[RA_Mul.scala 446:9:@4551.4]
  assign Reduction_2_io_matrix_i_3_23 = Reduction_1_io_matrix_3_23; // @[RA_Mul.scala 446:9:@4552.4]
  assign Reduction_2_io_matrix_i_3_24 = Reduction_1_io_matrix_3_24; // @[RA_Mul.scala 446:9:@4553.4]
  assign Reduction_2_io_matrix_i_4_9 = Reduction_1_io_matrix_4_9; // @[RA_Mul.scala 446:9:@4570.4]
  assign Reduction_2_io_matrix_i_4_12 = Reduction_1_io_matrix_4_12; // @[RA_Mul.scala 446:9:@4573.4]
  assign Reduction_2_io_matrix_i_4_13 = Reduction_1_io_matrix_4_13; // @[RA_Mul.scala 446:9:@4574.4]
  assign Reduction_2_io_matrix_i_4_14 = Reduction_1_io_matrix_4_14; // @[RA_Mul.scala 446:9:@4575.4]
  assign Reduction_2_io_matrix_i_4_15 = Reduction_1_io_matrix_4_15; // @[RA_Mul.scala 446:9:@4576.4]
  assign Reduction_2_io_matrix_i_4_16 = Reduction_1_io_matrix_4_16; // @[RA_Mul.scala 446:9:@4577.4]
  assign Reduction_2_io_matrix_i_4_17 = Reduction_1_io_matrix_4_17; // @[RA_Mul.scala 446:9:@4578.4]
  assign Reduction_2_io_matrix_i_4_18 = Reduction_1_io_matrix_4_18; // @[RA_Mul.scala 446:9:@4579.4]
  assign Reduction_2_io_matrix_i_4_19 = Reduction_1_io_matrix_4_19; // @[RA_Mul.scala 446:9:@4580.4]
  assign Reduction_2_io_matrix_i_4_20 = Reduction_1_io_matrix_4_20; // @[RA_Mul.scala 446:9:@4581.4]
  assign Reduction_2_io_matrix_i_4_23 = Reduction_1_io_matrix_4_23; // @[RA_Mul.scala 446:9:@4584.4]
  assign Reduction_2_io_matrix_i_5_12 = Reduction_1_io_matrix_5_12; // @[RA_Mul.scala 446:9:@4605.4]
  assign Reduction_2_io_matrix_i_5_15 = Reduction_1_io_matrix_5_15; // @[RA_Mul.scala 446:9:@4608.4]
  assign Reduction_2_io_matrix_i_5_16 = Reduction_1_io_matrix_5_16; // @[RA_Mul.scala 446:9:@4609.4]
  assign Reduction_2_io_matrix_i_5_17 = Reduction_1_io_matrix_5_17; // @[RA_Mul.scala 446:9:@4610.4]
  assign Reduction_2_io_matrix_i_5_18 = Reduction_1_io_matrix_5_18; // @[RA_Mul.scala 446:9:@4611.4]
  assign Reduction_2_io_matrix_i_5_19 = Reduction_1_io_matrix_5_19; // @[RA_Mul.scala 446:9:@4612.4]
  assign Reduction_3_io_matrix_i_0_0 = Reduction_2_io_matrix_o_0_0; // @[RA_Mul.scala 537:9:@4756.4]
  assign Reduction_3_io_matrix_i_0_1 = Reduction_2_io_matrix_o_0_1; // @[RA_Mul.scala 537:9:@4757.4]
  assign Reduction_3_io_matrix_i_0_2 = Reduction_2_io_matrix_o_0_2; // @[RA_Mul.scala 537:9:@4758.4]
  assign Reduction_3_io_matrix_i_0_3 = Reduction_2_io_matrix_o_0_3; // @[RA_Mul.scala 537:9:@4759.4]
  assign Reduction_3_io_matrix_i_0_4 = Reduction_2_io_matrix_o_0_4; // @[RA_Mul.scala 537:9:@4760.4]
  assign Reduction_3_io_matrix_i_0_5 = Reduction_2_io_matrix_o_0_5; // @[RA_Mul.scala 537:9:@4761.4]
  assign Reduction_3_io_matrix_i_0_6 = Reduction_2_io_matrix_o_0_6; // @[RA_Mul.scala 537:9:@4762.4]
  assign Reduction_3_io_matrix_i_0_7 = Reduction_2_io_matrix_o_0_7; // @[RA_Mul.scala 537:9:@4763.4]
  assign Reduction_3_io_matrix_i_0_8 = Reduction_2_io_matrix_o_0_8; // @[RA_Mul.scala 537:9:@4764.4]
  assign Reduction_3_io_matrix_i_0_9 = Reduction_2_io_matrix_o_0_9; // @[RA_Mul.scala 537:9:@4765.4]
  assign Reduction_3_io_matrix_i_0_10 = Reduction_2_io_matrix_o_0_10; // @[RA_Mul.scala 537:9:@4766.4]
  assign Reduction_3_io_matrix_i_0_11 = Reduction_2_io_matrix_o_0_11; // @[RA_Mul.scala 537:9:@4767.4]
  assign Reduction_3_io_matrix_i_0_12 = Reduction_2_io_matrix_o_0_12; // @[RA_Mul.scala 537:9:@4768.4]
  assign Reduction_3_io_matrix_i_0_13 = Reduction_2_io_matrix_o_0_13; // @[RA_Mul.scala 537:9:@4769.4]
  assign Reduction_3_io_matrix_i_0_14 = Reduction_2_io_matrix_o_0_14; // @[RA_Mul.scala 537:9:@4770.4]
  assign Reduction_3_io_matrix_i_0_15 = Reduction_2_io_matrix_o_0_15; // @[RA_Mul.scala 537:9:@4771.4]
  assign Reduction_3_io_matrix_i_0_16 = Reduction_2_io_matrix_o_0_16; // @[RA_Mul.scala 537:9:@4772.4]
  assign Reduction_3_io_matrix_i_0_17 = Reduction_2_io_matrix_o_0_17; // @[RA_Mul.scala 537:9:@4773.4]
  assign Reduction_3_io_matrix_i_0_18 = Reduction_2_io_matrix_o_0_18; // @[RA_Mul.scala 537:9:@4774.4]
  assign Reduction_3_io_matrix_i_0_19 = Reduction_2_io_matrix_o_0_19; // @[RA_Mul.scala 537:9:@4775.4]
  assign Reduction_3_io_matrix_i_0_20 = Reduction_2_io_matrix_o_0_20; // @[RA_Mul.scala 537:9:@4776.4]
  assign Reduction_3_io_matrix_i_0_21 = Reduction_2_io_matrix_o_0_21; // @[RA_Mul.scala 537:9:@4777.4]
  assign Reduction_3_io_matrix_i_0_22 = Reduction_2_io_matrix_o_0_22; // @[RA_Mul.scala 537:9:@4778.4]
  assign Reduction_3_io_matrix_i_0_23 = Reduction_2_io_matrix_o_0_23; // @[RA_Mul.scala 537:9:@4779.4]
  assign Reduction_3_io_matrix_i_0_24 = Reduction_2_io_matrix_o_0_24; // @[RA_Mul.scala 537:9:@4780.4]
  assign Reduction_3_io_matrix_i_0_25 = Reduction_2_io_matrix_o_0_25; // @[RA_Mul.scala 537:9:@4781.4]
  assign Reduction_3_io_matrix_i_0_26 = Reduction_2_io_matrix_o_0_26; // @[RA_Mul.scala 537:9:@4782.4]
  assign Reduction_3_io_matrix_i_0_27 = Reduction_2_io_matrix_o_0_27; // @[RA_Mul.scala 537:9:@4783.4]
  assign Reduction_3_io_matrix_i_0_28 = Reduction_2_io_matrix_o_0_28; // @[RA_Mul.scala 537:9:@4784.4]
  assign Reduction_3_io_matrix_i_0_29 = Reduction_2_io_matrix_o_0_29; // @[RA_Mul.scala 537:9:@4785.4]
  assign Reduction_3_io_matrix_i_0_30 = Reduction_2_io_matrix_o_0_30; // @[RA_Mul.scala 537:9:@4786.4]
  assign Reduction_3_io_matrix_i_0_31 = Reduction_2_io_matrix_o_0_31; // @[RA_Mul.scala 537:9:@4787.4]
  assign Reduction_3_io_matrix_i_1_2 = Reduction_2_io_matrix_o_1_2; // @[RA_Mul.scala 537:9:@4790.4]
  assign Reduction_3_io_matrix_i_1_4 = Reduction_2_io_matrix_o_1_4; // @[RA_Mul.scala 537:9:@4792.4]
  assign Reduction_3_io_matrix_i_1_5 = Reduction_2_io_matrix_o_1_5; // @[RA_Mul.scala 537:9:@4793.4]
  assign Reduction_3_io_matrix_i_1_6 = Reduction_2_io_matrix_o_1_6; // @[RA_Mul.scala 537:9:@4794.4]
  assign Reduction_3_io_matrix_i_1_7 = Reduction_2_io_matrix_o_1_7; // @[RA_Mul.scala 537:9:@4795.4]
  assign Reduction_3_io_matrix_i_1_8 = Reduction_2_io_matrix_o_1_8; // @[RA_Mul.scala 537:9:@4796.4]
  assign Reduction_3_io_matrix_i_1_9 = Reduction_2_io_matrix_o_1_9; // @[RA_Mul.scala 537:9:@4797.4]
  assign Reduction_3_io_matrix_i_1_10 = Reduction_2_io_matrix_o_1_10; // @[RA_Mul.scala 537:9:@4798.4]
  assign Reduction_3_io_matrix_i_1_11 = Reduction_2_io_matrix_o_1_11; // @[RA_Mul.scala 537:9:@4799.4]
  assign Reduction_3_io_matrix_i_1_12 = Reduction_2_io_matrix_o_1_12; // @[RA_Mul.scala 537:9:@4800.4]
  assign Reduction_3_io_matrix_i_1_13 = Reduction_2_io_matrix_o_1_13; // @[RA_Mul.scala 537:9:@4801.4]
  assign Reduction_3_io_matrix_i_1_14 = Reduction_2_io_matrix_o_1_14; // @[RA_Mul.scala 537:9:@4802.4]
  assign Reduction_3_io_matrix_i_1_15 = Reduction_2_io_matrix_o_1_15; // @[RA_Mul.scala 537:9:@4803.4]
  assign Reduction_3_io_matrix_i_1_16 = Reduction_2_io_matrix_o_1_16; // @[RA_Mul.scala 537:9:@4804.4]
  assign Reduction_3_io_matrix_i_1_17 = Reduction_2_io_matrix_o_1_17; // @[RA_Mul.scala 537:9:@4805.4]
  assign Reduction_3_io_matrix_i_1_18 = Reduction_2_io_matrix_o_1_18; // @[RA_Mul.scala 537:9:@4806.4]
  assign Reduction_3_io_matrix_i_1_19 = Reduction_2_io_matrix_o_1_19; // @[RA_Mul.scala 537:9:@4807.4]
  assign Reduction_3_io_matrix_i_1_20 = Reduction_2_io_matrix_o_1_20; // @[RA_Mul.scala 537:9:@4808.4]
  assign Reduction_3_io_matrix_i_1_21 = Reduction_2_io_matrix_o_1_21; // @[RA_Mul.scala 537:9:@4809.4]
  assign Reduction_3_io_matrix_i_1_22 = Reduction_2_io_matrix_o_1_22; // @[RA_Mul.scala 537:9:@4810.4]
  assign Reduction_3_io_matrix_i_1_23 = Reduction_2_io_matrix_o_1_23; // @[RA_Mul.scala 537:9:@4811.4]
  assign Reduction_3_io_matrix_i_1_24 = Reduction_2_io_matrix_o_1_24; // @[RA_Mul.scala 537:9:@4812.4]
  assign Reduction_3_io_matrix_i_1_25 = Reduction_2_io_matrix_o_1_25; // @[RA_Mul.scala 537:9:@4813.4]
  assign Reduction_3_io_matrix_i_1_26 = Reduction_2_io_matrix_o_1_26; // @[RA_Mul.scala 537:9:@4814.4]
  assign Reduction_3_io_matrix_i_1_27 = Reduction_2_io_matrix_o_1_27; // @[RA_Mul.scala 537:9:@4815.4]
  assign Reduction_3_io_matrix_i_1_28 = Reduction_2_io_matrix_o_1_28; // @[RA_Mul.scala 537:9:@4816.4]
  assign Reduction_3_io_matrix_i_1_30 = Reduction_2_io_matrix_o_1_30; // @[RA_Mul.scala 537:9:@4818.4]
  assign Reduction_3_io_matrix_i_2_4 = Reduction_2_io_matrix_o_2_4; // @[RA_Mul.scala 537:9:@4824.4]
  assign Reduction_3_io_matrix_i_2_9 = Reduction_2_io_matrix_o_2_9; // @[RA_Mul.scala 537:9:@4829.4]
  assign Reduction_3_io_matrix_i_2_10 = Reduction_2_io_matrix_o_2_10; // @[RA_Mul.scala 537:9:@4830.4]
  assign Reduction_3_io_matrix_i_2_11 = Reduction_2_io_matrix_o_2_11; // @[RA_Mul.scala 537:9:@4831.4]
  assign Reduction_3_io_matrix_i_2_12 = Reduction_2_io_matrix_o_2_12; // @[RA_Mul.scala 537:9:@4832.4]
  assign Reduction_3_io_matrix_i_2_13 = Reduction_2_io_matrix_o_2_13; // @[RA_Mul.scala 537:9:@4833.4]
  assign Reduction_3_io_matrix_i_2_14 = Reduction_2_io_matrix_o_2_14; // @[RA_Mul.scala 537:9:@4834.4]
  assign Reduction_3_io_matrix_i_2_15 = Reduction_2_io_matrix_o_2_15; // @[RA_Mul.scala 537:9:@4835.4]
  assign Reduction_3_io_matrix_i_2_16 = Reduction_2_io_matrix_o_2_16; // @[RA_Mul.scala 537:9:@4836.4]
  assign Reduction_3_io_matrix_i_2_17 = Reduction_2_io_matrix_o_2_17; // @[RA_Mul.scala 537:9:@4837.4]
  assign Reduction_3_io_matrix_i_2_18 = Reduction_2_io_matrix_o_2_18; // @[RA_Mul.scala 537:9:@4838.4]
  assign Reduction_3_io_matrix_i_2_19 = Reduction_2_io_matrix_o_2_19; // @[RA_Mul.scala 537:9:@4839.4]
  assign Reduction_3_io_matrix_i_2_20 = Reduction_2_io_matrix_o_2_20; // @[RA_Mul.scala 537:9:@4840.4]
  assign Reduction_3_io_matrix_i_2_21 = Reduction_2_io_matrix_o_2_21; // @[RA_Mul.scala 537:9:@4841.4]
  assign Reduction_3_io_matrix_i_2_22 = Reduction_2_io_matrix_o_2_22; // @[RA_Mul.scala 537:9:@4842.4]
  assign Reduction_3_io_matrix_i_2_23 = Reduction_2_io_matrix_o_2_23; // @[RA_Mul.scala 537:9:@4843.4]
  assign Reduction_3_io_matrix_i_2_24 = Reduction_2_io_matrix_o_2_24; // @[RA_Mul.scala 537:9:@4844.4]
  assign Reduction_3_io_matrix_i_2_27 = Reduction_2_io_matrix_o_2_27; // @[RA_Mul.scala 537:9:@4847.4]
  assign Reduction_3_io_matrix_i_2_30 = Reduction_2_io_matrix_o_2_30; // @[RA_Mul.scala 537:9:@4850.4]
  assign Reduction_3_io_matrix_i_3_9 = Reduction_2_io_matrix_o_3_9; // @[RA_Mul.scala 537:9:@4861.4]
  assign Reduction_3_io_matrix_i_3_13 = Reduction_2_io_matrix_o_3_13; // @[RA_Mul.scala 537:9:@4865.4]
  assign Reduction_3_io_matrix_i_3_14 = Reduction_2_io_matrix_o_3_14; // @[RA_Mul.scala 537:9:@4866.4]
  assign Reduction_3_io_matrix_i_3_15 = Reduction_2_io_matrix_o_3_15; // @[RA_Mul.scala 537:9:@4867.4]
  assign Reduction_3_io_matrix_i_3_16 = Reduction_2_io_matrix_o_3_16; // @[RA_Mul.scala 537:9:@4868.4]
  assign Reduction_3_io_matrix_i_3_17 = Reduction_2_io_matrix_o_3_17; // @[RA_Mul.scala 537:9:@4869.4]
  assign Reduction_3_io_matrix_i_3_18 = Reduction_2_io_matrix_o_3_18; // @[RA_Mul.scala 537:9:@4870.4]
  assign Reduction_3_io_matrix_i_3_19 = Reduction_2_io_matrix_o_3_19; // @[RA_Mul.scala 537:9:@4871.4]
  assign Reduction_3_io_matrix_i_3_20 = Reduction_2_io_matrix_o_3_20; // @[RA_Mul.scala 537:9:@4872.4]
  assign Reduction_3_io_matrix_i_3_21 = Reduction_2_io_matrix_o_3_21; // @[RA_Mul.scala 537:9:@4873.4]
  assign Reduction_3_io_matrix_i_3_23 = Reduction_2_io_matrix_o_3_23; // @[RA_Mul.scala 537:9:@4875.4]
  assign Reduction_4_io_matrix_i_0_0 = Reduction_3_io_matrix_o_0_0; // @[RA_Mul.scala 600:9:@4983.4]
  assign Reduction_4_io_matrix_i_0_1 = Reduction_3_io_matrix_o_0_1; // @[RA_Mul.scala 600:9:@4984.4]
  assign Reduction_4_io_matrix_i_0_2 = Reduction_3_io_matrix_o_0_2; // @[RA_Mul.scala 600:9:@4985.4]
  assign Reduction_4_io_matrix_i_0_3 = Reduction_3_io_matrix_o_0_3; // @[RA_Mul.scala 600:9:@4986.4]
  assign Reduction_4_io_matrix_i_0_4 = Reduction_3_io_matrix_o_0_4; // @[RA_Mul.scala 600:9:@4987.4]
  assign Reduction_4_io_matrix_i_0_5 = Reduction_3_io_matrix_o_0_5; // @[RA_Mul.scala 600:9:@4988.4]
  assign Reduction_4_io_matrix_i_0_6 = Reduction_3_io_matrix_o_0_6; // @[RA_Mul.scala 600:9:@4989.4]
  assign Reduction_4_io_matrix_i_0_7 = Reduction_3_io_matrix_o_0_7; // @[RA_Mul.scala 600:9:@4990.4]
  assign Reduction_4_io_matrix_i_0_8 = Reduction_3_io_matrix_o_0_8; // @[RA_Mul.scala 600:9:@4991.4]
  assign Reduction_4_io_matrix_i_0_9 = Reduction_3_io_matrix_o_0_9; // @[RA_Mul.scala 600:9:@4992.4]
  assign Reduction_4_io_matrix_i_0_10 = Reduction_3_io_matrix_o_0_10; // @[RA_Mul.scala 600:9:@4993.4]
  assign Reduction_4_io_matrix_i_0_11 = Reduction_3_io_matrix_o_0_11; // @[RA_Mul.scala 600:9:@4994.4]
  assign Reduction_4_io_matrix_i_0_12 = Reduction_3_io_matrix_o_0_12; // @[RA_Mul.scala 600:9:@4995.4]
  assign Reduction_4_io_matrix_i_0_13 = Reduction_3_io_matrix_o_0_13; // @[RA_Mul.scala 600:9:@4996.4]
  assign Reduction_4_io_matrix_i_0_14 = Reduction_3_io_matrix_o_0_14; // @[RA_Mul.scala 600:9:@4997.4]
  assign Reduction_4_io_matrix_i_0_15 = Reduction_3_io_matrix_o_0_15; // @[RA_Mul.scala 600:9:@4998.4]
  assign Reduction_4_io_matrix_i_0_16 = Reduction_3_io_matrix_o_0_16; // @[RA_Mul.scala 600:9:@4999.4]
  assign Reduction_4_io_matrix_i_0_17 = Reduction_3_io_matrix_o_0_17; // @[RA_Mul.scala 600:9:@5000.4]
  assign Reduction_4_io_matrix_i_0_18 = Reduction_3_io_matrix_o_0_18; // @[RA_Mul.scala 600:9:@5001.4]
  assign Reduction_4_io_matrix_i_0_19 = Reduction_3_io_matrix_o_0_19; // @[RA_Mul.scala 600:9:@5002.4]
  assign Reduction_4_io_matrix_i_0_20 = Reduction_3_io_matrix_o_0_20; // @[RA_Mul.scala 600:9:@5003.4]
  assign Reduction_4_io_matrix_i_0_21 = Reduction_3_io_matrix_o_0_21; // @[RA_Mul.scala 600:9:@5004.4]
  assign Reduction_4_io_matrix_i_0_22 = Reduction_3_io_matrix_o_0_22; // @[RA_Mul.scala 600:9:@5005.4]
  assign Reduction_4_io_matrix_i_0_23 = Reduction_3_io_matrix_o_0_23; // @[RA_Mul.scala 600:9:@5006.4]
  assign Reduction_4_io_matrix_i_0_24 = Reduction_3_io_matrix_o_0_24; // @[RA_Mul.scala 600:9:@5007.4]
  assign Reduction_4_io_matrix_i_0_25 = Reduction_3_io_matrix_o_0_25; // @[RA_Mul.scala 600:9:@5008.4]
  assign Reduction_4_io_matrix_i_0_26 = Reduction_3_io_matrix_o_0_26; // @[RA_Mul.scala 600:9:@5009.4]
  assign Reduction_4_io_matrix_i_0_27 = Reduction_3_io_matrix_o_0_27; // @[RA_Mul.scala 600:9:@5010.4]
  assign Reduction_4_io_matrix_i_0_28 = Reduction_3_io_matrix_o_0_28; // @[RA_Mul.scala 600:9:@5011.4]
  assign Reduction_4_io_matrix_i_0_29 = Reduction_3_io_matrix_o_0_29; // @[RA_Mul.scala 600:9:@5012.4]
  assign Reduction_4_io_matrix_i_0_30 = Reduction_3_io_matrix_o_0_30; // @[RA_Mul.scala 600:9:@5013.4]
  assign Reduction_4_io_matrix_i_0_31 = Reduction_3_io_matrix_o_0_31; // @[RA_Mul.scala 600:9:@5014.4]
  assign Reduction_4_io_matrix_i_1_3 = Reduction_3_io_matrix_o_1_3; // @[RA_Mul.scala 600:9:@5018.4]
  assign Reduction_4_io_matrix_i_1_5 = Reduction_3_io_matrix_o_1_5; // @[RA_Mul.scala 600:9:@5020.4]
  assign Reduction_4_io_matrix_i_1_6 = Reduction_3_io_matrix_o_1_6; // @[RA_Mul.scala 600:9:@5021.4]
  assign Reduction_4_io_matrix_i_1_7 = Reduction_3_io_matrix_o_1_7; // @[RA_Mul.scala 600:9:@5022.4]
  assign Reduction_4_io_matrix_i_1_8 = Reduction_3_io_matrix_o_1_8; // @[RA_Mul.scala 600:9:@5023.4]
  assign Reduction_4_io_matrix_i_1_9 = Reduction_3_io_matrix_o_1_9; // @[RA_Mul.scala 600:9:@5024.4]
  assign Reduction_4_io_matrix_i_1_10 = Reduction_3_io_matrix_o_1_10; // @[RA_Mul.scala 600:9:@5025.4]
  assign Reduction_4_io_matrix_i_1_11 = Reduction_3_io_matrix_o_1_11; // @[RA_Mul.scala 600:9:@5026.4]
  assign Reduction_4_io_matrix_i_1_12 = Reduction_3_io_matrix_o_1_12; // @[RA_Mul.scala 600:9:@5027.4]
  assign Reduction_4_io_matrix_i_1_13 = Reduction_3_io_matrix_o_1_13; // @[RA_Mul.scala 600:9:@5028.4]
  assign Reduction_4_io_matrix_i_1_14 = Reduction_3_io_matrix_o_1_14; // @[RA_Mul.scala 600:9:@5029.4]
  assign Reduction_4_io_matrix_i_1_15 = Reduction_3_io_matrix_o_1_15; // @[RA_Mul.scala 600:9:@5030.4]
  assign Reduction_4_io_matrix_i_1_16 = Reduction_3_io_matrix_o_1_16; // @[RA_Mul.scala 600:9:@5031.4]
  assign Reduction_4_io_matrix_i_1_17 = Reduction_3_io_matrix_o_1_17; // @[RA_Mul.scala 600:9:@5032.4]
  assign Reduction_4_io_matrix_i_1_18 = Reduction_3_io_matrix_o_1_18; // @[RA_Mul.scala 600:9:@5033.4]
  assign Reduction_4_io_matrix_i_1_19 = Reduction_3_io_matrix_o_1_19; // @[RA_Mul.scala 600:9:@5034.4]
  assign Reduction_4_io_matrix_i_1_20 = Reduction_3_io_matrix_o_1_20; // @[RA_Mul.scala 600:9:@5035.4]
  assign Reduction_4_io_matrix_i_1_21 = Reduction_3_io_matrix_o_1_21; // @[RA_Mul.scala 600:9:@5036.4]
  assign Reduction_4_io_matrix_i_1_22 = Reduction_3_io_matrix_o_1_22; // @[RA_Mul.scala 600:9:@5037.4]
  assign Reduction_4_io_matrix_i_1_23 = Reduction_3_io_matrix_o_1_23; // @[RA_Mul.scala 600:9:@5038.4]
  assign Reduction_4_io_matrix_i_1_24 = Reduction_3_io_matrix_o_1_24; // @[RA_Mul.scala 600:9:@5039.4]
  assign Reduction_4_io_matrix_i_1_25 = Reduction_3_io_matrix_o_1_25; // @[RA_Mul.scala 600:9:@5040.4]
  assign Reduction_4_io_matrix_i_1_26 = Reduction_3_io_matrix_o_1_26; // @[RA_Mul.scala 600:9:@5041.4]
  assign Reduction_4_io_matrix_i_1_28 = Reduction_3_io_matrix_o_1_28; // @[RA_Mul.scala 600:9:@5043.4]
  assign Reduction_4_io_matrix_i_1_31 = Reduction_3_io_matrix_o_1_31; // @[RA_Mul.scala 600:9:@5046.4]
  assign Reduction_4_io_matrix_i_2_5 = Reduction_3_io_matrix_o_2_5; // @[RA_Mul.scala 600:9:@5052.4]
  assign Reduction_4_io_matrix_i_2_13 = Reduction_3_io_matrix_o_2_13; // @[RA_Mul.scala 600:9:@5060.4]
  assign Reduction_4_io_matrix_i_2_14 = Reduction_3_io_matrix_o_2_14; // @[RA_Mul.scala 600:9:@5061.4]
  assign Reduction_4_io_matrix_i_2_15 = Reduction_3_io_matrix_o_2_15; // @[RA_Mul.scala 600:9:@5062.4]
  assign Reduction_4_io_matrix_i_2_16 = Reduction_3_io_matrix_o_2_16; // @[RA_Mul.scala 600:9:@5063.4]
  assign Reduction_4_io_matrix_i_2_17 = Reduction_3_io_matrix_o_2_17; // @[RA_Mul.scala 600:9:@5064.4]
  assign Reduction_4_io_matrix_i_2_18 = Reduction_3_io_matrix_o_2_18; // @[RA_Mul.scala 600:9:@5065.4]
  assign Reduction_4_io_matrix_i_2_19 = Reduction_3_io_matrix_o_2_19; // @[RA_Mul.scala 600:9:@5066.4]
  assign Reduction_4_io_matrix_i_2_20 = Reduction_3_io_matrix_o_2_20; // @[RA_Mul.scala 600:9:@5067.4]
  assign Reduction_4_io_matrix_i_2_21 = Reduction_3_io_matrix_o_2_21; // @[RA_Mul.scala 600:9:@5068.4]
  assign Reduction_4_io_matrix_i_2_23 = Reduction_3_io_matrix_o_2_23; // @[RA_Mul.scala 600:9:@5070.4]
  assign Reduction_4_io_matrix_i_2_25 = Reduction_3_io_matrix_o_2_25; // @[RA_Mul.scala 600:9:@5072.4]
  assign Reduction_4_io_matrix_i_2_28 = Reduction_3_io_matrix_o_2_28; // @[RA_Mul.scala 600:9:@5075.4]
  assign PPLRegs2_clock = clock; // @[:@5144.4]
  assign PPLRegs2_reset = reset; // @[:@5145.4]
  assign PPLRegs2_io_matrix_i_0_0 = Reduction_4_io_matrix_o_0_0; // @[RA_Mul.scala 715:9:@5210.4]
  assign PPLRegs2_io_matrix_i_0_1 = Reduction_4_io_matrix_o_0_1; // @[RA_Mul.scala 715:9:@5211.4]
  assign PPLRegs2_io_matrix_i_0_2 = Reduction_4_io_matrix_o_0_2; // @[RA_Mul.scala 715:9:@5212.4]
  assign PPLRegs2_io_matrix_i_0_3 = Reduction_4_io_matrix_o_0_3; // @[RA_Mul.scala 715:9:@5213.4]
  assign PPLRegs2_io_matrix_i_0_4 = Reduction_4_io_matrix_o_0_4; // @[RA_Mul.scala 715:9:@5214.4]
  assign PPLRegs2_io_matrix_i_0_5 = Reduction_4_io_matrix_o_0_5; // @[RA_Mul.scala 715:9:@5215.4]
  assign PPLRegs2_io_matrix_i_0_6 = Reduction_4_io_matrix_o_0_6; // @[RA_Mul.scala 715:9:@5216.4]
  assign PPLRegs2_io_matrix_i_0_7 = Reduction_4_io_matrix_o_0_7; // @[RA_Mul.scala 715:9:@5217.4]
  assign PPLRegs2_io_matrix_i_0_8 = Reduction_4_io_matrix_o_0_8; // @[RA_Mul.scala 715:9:@5218.4]
  assign PPLRegs2_io_matrix_i_0_9 = Reduction_4_io_matrix_o_0_9; // @[RA_Mul.scala 715:9:@5219.4]
  assign PPLRegs2_io_matrix_i_0_10 = Reduction_4_io_matrix_o_0_10; // @[RA_Mul.scala 715:9:@5220.4]
  assign PPLRegs2_io_matrix_i_0_11 = Reduction_4_io_matrix_o_0_11; // @[RA_Mul.scala 715:9:@5221.4]
  assign PPLRegs2_io_matrix_i_0_12 = Reduction_4_io_matrix_o_0_12; // @[RA_Mul.scala 715:9:@5222.4]
  assign PPLRegs2_io_matrix_i_0_13 = Reduction_4_io_matrix_o_0_13; // @[RA_Mul.scala 715:9:@5223.4]
  assign PPLRegs2_io_matrix_i_0_14 = Reduction_4_io_matrix_o_0_14; // @[RA_Mul.scala 715:9:@5224.4]
  assign PPLRegs2_io_matrix_i_0_15 = Reduction_4_io_matrix_o_0_15; // @[RA_Mul.scala 715:9:@5225.4]
  assign PPLRegs2_io_matrix_i_0_16 = Reduction_4_io_matrix_o_0_16; // @[RA_Mul.scala 715:9:@5226.4]
  assign PPLRegs2_io_matrix_i_0_17 = Reduction_4_io_matrix_o_0_17; // @[RA_Mul.scala 715:9:@5227.4]
  assign PPLRegs2_io_matrix_i_0_18 = Reduction_4_io_matrix_o_0_18; // @[RA_Mul.scala 715:9:@5228.4]
  assign PPLRegs2_io_matrix_i_0_19 = Reduction_4_io_matrix_o_0_19; // @[RA_Mul.scala 715:9:@5229.4]
  assign PPLRegs2_io_matrix_i_0_20 = Reduction_4_io_matrix_o_0_20; // @[RA_Mul.scala 715:9:@5230.4]
  assign PPLRegs2_io_matrix_i_0_21 = Reduction_4_io_matrix_o_0_21; // @[RA_Mul.scala 715:9:@5231.4]
  assign PPLRegs2_io_matrix_i_0_22 = Reduction_4_io_matrix_o_0_22; // @[RA_Mul.scala 715:9:@5232.4]
  assign PPLRegs2_io_matrix_i_0_23 = Reduction_4_io_matrix_o_0_23; // @[RA_Mul.scala 715:9:@5233.4]
  assign PPLRegs2_io_matrix_i_0_24 = Reduction_4_io_matrix_o_0_24; // @[RA_Mul.scala 715:9:@5234.4]
  assign PPLRegs2_io_matrix_i_0_25 = Reduction_4_io_matrix_o_0_25; // @[RA_Mul.scala 715:9:@5235.4]
  assign PPLRegs2_io_matrix_i_0_26 = Reduction_4_io_matrix_o_0_26; // @[RA_Mul.scala 715:9:@5236.4]
  assign PPLRegs2_io_matrix_i_0_27 = Reduction_4_io_matrix_o_0_27; // @[RA_Mul.scala 715:9:@5237.4]
  assign PPLRegs2_io_matrix_i_0_28 = Reduction_4_io_matrix_o_0_28; // @[RA_Mul.scala 715:9:@5238.4]
  assign PPLRegs2_io_matrix_i_0_29 = Reduction_4_io_matrix_o_0_29; // @[RA_Mul.scala 715:9:@5239.4]
  assign PPLRegs2_io_matrix_i_0_30 = Reduction_4_io_matrix_o_0_30; // @[RA_Mul.scala 715:9:@5240.4]
  assign PPLRegs2_io_matrix_i_0_31 = Reduction_4_io_matrix_o_0_31; // @[RA_Mul.scala 715:9:@5241.4]
  assign PPLRegs2_io_matrix_i_1_4 = Reduction_4_io_matrix_o_1_4; // @[RA_Mul.scala 715:9:@5246.4]
  assign PPLRegs2_io_matrix_i_1_6 = Reduction_4_io_matrix_o_1_6; // @[RA_Mul.scala 715:9:@5248.4]
  assign PPLRegs2_io_matrix_i_1_7 = Reduction_4_io_matrix_o_1_7; // @[RA_Mul.scala 715:9:@5249.4]
  assign PPLRegs2_io_matrix_i_1_8 = Reduction_4_io_matrix_o_1_8; // @[RA_Mul.scala 715:9:@5250.4]
  assign PPLRegs2_io_matrix_i_1_9 = Reduction_4_io_matrix_o_1_9; // @[RA_Mul.scala 715:9:@5251.4]
  assign PPLRegs2_io_matrix_i_1_10 = Reduction_4_io_matrix_o_1_10; // @[RA_Mul.scala 715:9:@5252.4]
  assign PPLRegs2_io_matrix_i_1_11 = Reduction_4_io_matrix_o_1_11; // @[RA_Mul.scala 715:9:@5253.4]
  assign PPLRegs2_io_matrix_i_1_12 = Reduction_4_io_matrix_o_1_12; // @[RA_Mul.scala 715:9:@5254.4]
  assign PPLRegs2_io_matrix_i_1_13 = Reduction_4_io_matrix_o_1_13; // @[RA_Mul.scala 715:9:@5255.4]
  assign PPLRegs2_io_matrix_i_1_14 = Reduction_4_io_matrix_o_1_14; // @[RA_Mul.scala 715:9:@5256.4]
  assign PPLRegs2_io_matrix_i_1_15 = Reduction_4_io_matrix_o_1_15; // @[RA_Mul.scala 715:9:@5257.4]
  assign PPLRegs2_io_matrix_i_1_16 = Reduction_4_io_matrix_o_1_16; // @[RA_Mul.scala 715:9:@5258.4]
  assign PPLRegs2_io_matrix_i_1_17 = Reduction_4_io_matrix_o_1_17; // @[RA_Mul.scala 715:9:@5259.4]
  assign PPLRegs2_io_matrix_i_1_18 = Reduction_4_io_matrix_o_1_18; // @[RA_Mul.scala 715:9:@5260.4]
  assign PPLRegs2_io_matrix_i_1_19 = Reduction_4_io_matrix_o_1_19; // @[RA_Mul.scala 715:9:@5261.4]
  assign PPLRegs2_io_matrix_i_1_20 = Reduction_4_io_matrix_o_1_20; // @[RA_Mul.scala 715:9:@5262.4]
  assign PPLRegs2_io_matrix_i_1_21 = Reduction_4_io_matrix_o_1_21; // @[RA_Mul.scala 715:9:@5263.4]
  assign PPLRegs2_io_matrix_i_1_22 = Reduction_4_io_matrix_o_1_22; // @[RA_Mul.scala 715:9:@5264.4]
  assign PPLRegs2_io_matrix_i_1_23 = Reduction_4_io_matrix_o_1_23; // @[RA_Mul.scala 715:9:@5265.4]
  assign PPLRegs2_io_matrix_i_1_24 = Reduction_4_io_matrix_o_1_24; // @[RA_Mul.scala 715:9:@5266.4]
  assign PPLRegs2_io_matrix_i_1_25 = Reduction_4_io_matrix_o_1_25; // @[RA_Mul.scala 715:9:@5267.4]
  assign PPLRegs2_io_matrix_i_1_26 = Reduction_4_io_matrix_o_1_26; // @[RA_Mul.scala 715:9:@5268.4]
  assign PPLRegs2_io_matrix_i_1_27 = Reduction_4_io_matrix_o_1_27; // @[RA_Mul.scala 715:9:@5269.4]
  assign PPLRegs2_io_matrix_i_1_29 = Reduction_4_io_matrix_o_1_29; // @[RA_Mul.scala 715:9:@5271.4]
  assign PPLRegs2_io_matrix_i_1_31 = Reduction_4_io_matrix_o_1_31; // @[RA_Mul.scala 715:9:@5273.4]
  assign TailAdder_io_B = {_T_3139,_T_3124}; // @[RA_Mul.scala 619:14:@5340.4]
  assign TailAdder_io_A = {_T_3108,_T_3093}; // @[RA_Mul.scala 618:14:@5339.4]
  assign PPLRegs3_clock = clock; // @[:@5343.4]
  assign PPLRegs3_reset = reset; // @[:@5344.4]
  assign PPLRegs3_io_S_i = TailAdder_io_S; // @[RA_Mul.scala 730:16:@5345.4]
endmodule
