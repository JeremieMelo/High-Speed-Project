module PPGen( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [15:0] io_PP_0, // @[:@6.4]
  output [15:0] io_PP_1, // @[:@6.4]
  output [15:0] io_PP_2, // @[:@6.4]
  output [15:0] io_PP_3, // @[:@6.4]
  output [15:0] io_PP_4, // @[:@6.4]
  output [15:0] io_PP_5, // @[:@6.4]
  output [15:0] io_PP_6, // @[:@6.4]
  output [15:0] io_PP_7, // @[:@6.4]
  output [7:0]  io_SS, // @[:@6.4]
  output [7:0]  io_SC, // @[:@6.4]
  output [7:0]  io_S, // @[:@6.4]
  input  [2:0]  io_eB_0, // @[:@6.4]
  input  [2:0]  io_eB_1, // @[:@6.4]
  input  [2:0]  io_eB_2, // @[:@6.4]
  input  [2:0]  io_eB_3, // @[:@6.4]
  input  [2:0]  io_eB_4, // @[:@6.4]
  input  [2:0]  io_eB_5, // @[:@6.4]
  input  [2:0]  io_eB_6, // @[:@6.4]
  input  [2:0]  io_eB_7, // @[:@6.4]
  input  [15:0] io_A // @[:@6.4]
);
  wire  _T_93; // @[RA_Mul.scala 62:19:@11.4]
  wire  _T_95; // @[RA_Mul.scala 62:44:@12.4]
  wire  _T_96; // @[RA_Mul.scala 62:32:@13.4]
  wire  _T_99; // @[RA_Mul.scala 64:25:@18.6]
  wire  _T_101; // @[RA_Mul.scala 66:25:@23.8]
  wire [16:0] _GEN_40; // @[RA_Mul.scala 67:25:@25.10]
  wire [16:0] _T_102; // @[RA_Mul.scala 67:25:@25.10]
  wire [15:0] _T_103; // @[RA_Mul.scala 67:30:@26.10]
  wire  _T_105; // @[RA_Mul.scala 68:25:@30.10]
  wire [15:0] _T_106; // @[RA_Mul.scala 69:19:@32.12]
  wire  _T_108; // @[RA_Mul.scala 70:25:@36.12]
  wire [15:0] _T_111; // @[RA_Mul.scala 71:19:@40.14]
  wire [15:0] _GEN_0; // @[RA_Mul.scala 70:38:@37.12]
  wire [15:0] _GEN_1; // @[RA_Mul.scala 68:39:@31.10]
  wire [15:0] _GEN_2; // @[RA_Mul.scala 66:39:@24.8]
  wire [15:0] _GEN_3; // @[RA_Mul.scala 64:39:@19.6]
  wire  S_v_0; // @[RA_Mul.scala 76:23:@46.4]
  wire  _T_115; // @[RA_Mul.scala 77:36:@49.4]
  wire  _T_116; // @[RA_Mul.scala 77:30:@50.4]
  wire  SC_v_0; // @[RA_Mul.scala 77:16:@51.4]
  wire  _T_119; // @[RA_Mul.scala 62:19:@53.4]
  wire  _T_121; // @[RA_Mul.scala 62:44:@54.4]
  wire  _T_122; // @[RA_Mul.scala 62:32:@55.4]
  wire  _T_125; // @[RA_Mul.scala 64:25:@60.6]
  wire  _T_127; // @[RA_Mul.scala 66:25:@65.8]
  wire  _T_131; // @[RA_Mul.scala 68:25:@72.10]
  wire  _T_134; // @[RA_Mul.scala 70:25:@78.12]
  wire [15:0] _GEN_5; // @[RA_Mul.scala 70:38:@79.12]
  wire [15:0] _GEN_6; // @[RA_Mul.scala 68:39:@73.10]
  wire [15:0] _GEN_7; // @[RA_Mul.scala 66:39:@66.8]
  wire [15:0] _GEN_8; // @[RA_Mul.scala 64:39:@61.6]
  wire  S_v_1; // @[RA_Mul.scala 76:23:@88.4]
  wire  _T_142; // @[RA_Mul.scala 77:30:@92.4]
  wire  SC_v_1; // @[RA_Mul.scala 77:16:@93.4]
  wire  _T_145; // @[RA_Mul.scala 62:19:@95.4]
  wire  _T_147; // @[RA_Mul.scala 62:44:@96.4]
  wire  _T_148; // @[RA_Mul.scala 62:32:@97.4]
  wire  _T_151; // @[RA_Mul.scala 64:25:@102.6]
  wire  _T_153; // @[RA_Mul.scala 66:25:@107.8]
  wire  _T_157; // @[RA_Mul.scala 68:25:@114.10]
  wire  _T_160; // @[RA_Mul.scala 70:25:@120.12]
  wire [15:0] _GEN_10; // @[RA_Mul.scala 70:38:@121.12]
  wire [15:0] _GEN_11; // @[RA_Mul.scala 68:39:@115.10]
  wire [15:0] _GEN_12; // @[RA_Mul.scala 66:39:@108.8]
  wire [15:0] _GEN_13; // @[RA_Mul.scala 64:39:@103.6]
  wire  S_v_2; // @[RA_Mul.scala 76:23:@130.4]
  wire  _T_168; // @[RA_Mul.scala 77:30:@134.4]
  wire  SC_v_2; // @[RA_Mul.scala 77:16:@135.4]
  wire  _T_171; // @[RA_Mul.scala 62:19:@137.4]
  wire  _T_173; // @[RA_Mul.scala 62:44:@138.4]
  wire  _T_174; // @[RA_Mul.scala 62:32:@139.4]
  wire  _T_177; // @[RA_Mul.scala 64:25:@144.6]
  wire  _T_179; // @[RA_Mul.scala 66:25:@149.8]
  wire  _T_183; // @[RA_Mul.scala 68:25:@156.10]
  wire  _T_186; // @[RA_Mul.scala 70:25:@162.12]
  wire [15:0] _GEN_15; // @[RA_Mul.scala 70:38:@163.12]
  wire [15:0] _GEN_16; // @[RA_Mul.scala 68:39:@157.10]
  wire [15:0] _GEN_17; // @[RA_Mul.scala 66:39:@150.8]
  wire [15:0] _GEN_18; // @[RA_Mul.scala 64:39:@145.6]
  wire  S_v_3; // @[RA_Mul.scala 76:23:@172.4]
  wire  _T_194; // @[RA_Mul.scala 77:30:@176.4]
  wire  SC_v_3; // @[RA_Mul.scala 77:16:@177.4]
  wire  _T_197; // @[RA_Mul.scala 62:19:@179.4]
  wire  _T_199; // @[RA_Mul.scala 62:44:@180.4]
  wire  _T_200; // @[RA_Mul.scala 62:32:@181.4]
  wire  _T_203; // @[RA_Mul.scala 64:25:@186.6]
  wire  _T_205; // @[RA_Mul.scala 66:25:@191.8]
  wire  _T_209; // @[RA_Mul.scala 68:25:@198.10]
  wire  _T_212; // @[RA_Mul.scala 70:25:@204.12]
  wire [15:0] _GEN_20; // @[RA_Mul.scala 70:38:@205.12]
  wire [15:0] _GEN_21; // @[RA_Mul.scala 68:39:@199.10]
  wire [15:0] _GEN_22; // @[RA_Mul.scala 66:39:@192.8]
  wire [15:0] _GEN_23; // @[RA_Mul.scala 64:39:@187.6]
  wire  S_v_4; // @[RA_Mul.scala 76:23:@214.4]
  wire  _T_220; // @[RA_Mul.scala 77:30:@218.4]
  wire  SC_v_4; // @[RA_Mul.scala 77:16:@219.4]
  wire  _T_223; // @[RA_Mul.scala 62:19:@221.4]
  wire  _T_225; // @[RA_Mul.scala 62:44:@222.4]
  wire  _T_226; // @[RA_Mul.scala 62:32:@223.4]
  wire  _T_229; // @[RA_Mul.scala 64:25:@228.6]
  wire  _T_231; // @[RA_Mul.scala 66:25:@233.8]
  wire  _T_235; // @[RA_Mul.scala 68:25:@240.10]
  wire  _T_238; // @[RA_Mul.scala 70:25:@246.12]
  wire [15:0] _GEN_25; // @[RA_Mul.scala 70:38:@247.12]
  wire [15:0] _GEN_26; // @[RA_Mul.scala 68:39:@241.10]
  wire [15:0] _GEN_27; // @[RA_Mul.scala 66:39:@234.8]
  wire [15:0] _GEN_28; // @[RA_Mul.scala 64:39:@229.6]
  wire  S_v_5; // @[RA_Mul.scala 76:23:@256.4]
  wire  _T_246; // @[RA_Mul.scala 77:30:@260.4]
  wire  SC_v_5; // @[RA_Mul.scala 77:16:@261.4]
  wire  _T_249; // @[RA_Mul.scala 62:19:@263.4]
  wire  _T_251; // @[RA_Mul.scala 62:44:@264.4]
  wire  _T_252; // @[RA_Mul.scala 62:32:@265.4]
  wire  _T_255; // @[RA_Mul.scala 64:25:@270.6]
  wire  _T_257; // @[RA_Mul.scala 66:25:@275.8]
  wire  _T_261; // @[RA_Mul.scala 68:25:@282.10]
  wire  _T_264; // @[RA_Mul.scala 70:25:@288.12]
  wire [15:0] _GEN_30; // @[RA_Mul.scala 70:38:@289.12]
  wire [15:0] _GEN_31; // @[RA_Mul.scala 68:39:@283.10]
  wire [15:0] _GEN_32; // @[RA_Mul.scala 66:39:@276.8]
  wire [15:0] _GEN_33; // @[RA_Mul.scala 64:39:@271.6]
  wire  S_v_6; // @[RA_Mul.scala 76:23:@298.4]
  wire  _T_272; // @[RA_Mul.scala 77:30:@302.4]
  wire  SC_v_6; // @[RA_Mul.scala 77:16:@303.4]
  wire  _T_275; // @[RA_Mul.scala 62:19:@305.4]
  wire  _T_277; // @[RA_Mul.scala 62:44:@306.4]
  wire  _T_278; // @[RA_Mul.scala 62:32:@307.4]
  wire  _T_281; // @[RA_Mul.scala 64:25:@312.6]
  wire  _T_283; // @[RA_Mul.scala 66:25:@317.8]
  wire  _T_287; // @[RA_Mul.scala 68:25:@324.10]
  wire  _T_290; // @[RA_Mul.scala 70:25:@330.12]
  wire [15:0] _GEN_35; // @[RA_Mul.scala 70:38:@331.12]
  wire [15:0] _GEN_36; // @[RA_Mul.scala 68:39:@325.10]
  wire [15:0] _GEN_37; // @[RA_Mul.scala 66:39:@318.8]
  wire [15:0] _GEN_38; // @[RA_Mul.scala 64:39:@313.6]
  wire  S_v_7; // @[RA_Mul.scala 76:23:@340.4]
  wire  _T_298; // @[RA_Mul.scala 77:30:@344.4]
  wire  SC_v_7; // @[RA_Mul.scala 77:16:@345.4]
  wire [1:0] _T_300; // @[RA_Mul.scala 79:21:@347.4]
  wire [1:0] _T_301; // @[RA_Mul.scala 79:21:@348.4]
  wire [3:0] _T_302; // @[RA_Mul.scala 79:21:@349.4]
  wire [1:0] _T_303; // @[RA_Mul.scala 79:21:@350.4]
  wire [1:0] _T_304; // @[RA_Mul.scala 79:21:@351.4]
  wire [3:0] _T_305; // @[RA_Mul.scala 79:21:@352.4]
  wire [1:0] _T_307; // @[RA_Mul.scala 80:23:@355.4]
  wire [1:0] _T_308; // @[RA_Mul.scala 80:23:@356.4]
  wire [3:0] _T_309; // @[RA_Mul.scala 80:23:@357.4]
  wire [1:0] _T_310; // @[RA_Mul.scala 80:23:@358.4]
  wire [1:0] _T_311; // @[RA_Mul.scala 80:23:@359.4]
  wire [3:0] _T_312; // @[RA_Mul.scala 80:23:@360.4]
  assign _T_93 = io_eB_0 == 3'h0; // @[RA_Mul.scala 62:19:@11.4]
  assign _T_95 = io_eB_0 == 3'h4; // @[RA_Mul.scala 62:44:@12.4]
  assign _T_96 = _T_93 | _T_95; // @[RA_Mul.scala 62:32:@13.4]
  assign _T_99 = io_eB_0 == 3'h1; // @[RA_Mul.scala 64:25:@18.6]
  assign _T_101 = io_eB_0 == 3'h2; // @[RA_Mul.scala 66:25:@23.8]
  assign _GEN_40 = {{1'd0}, io_A}; // @[RA_Mul.scala 67:25:@25.10]
  assign _T_102 = _GEN_40 << 1; // @[RA_Mul.scala 67:25:@25.10]
  assign _T_103 = _T_102[15:0]; // @[RA_Mul.scala 67:30:@26.10]
  assign _T_105 = io_eB_0 == 3'h5; // @[RA_Mul.scala 68:25:@30.10]
  assign _T_106 = ~ io_A; // @[RA_Mul.scala 69:19:@32.12]
  assign _T_108 = io_eB_0 == 3'h6; // @[RA_Mul.scala 70:25:@36.12]
  assign _T_111 = ~ _T_103; // @[RA_Mul.scala 71:19:@40.14]
  assign _GEN_0 = _T_108 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@37.12]
  assign _GEN_1 = _T_105 ? _T_106 : _GEN_0; // @[RA_Mul.scala 68:39:@31.10]
  assign _GEN_2 = _T_101 ? _T_103 : _GEN_1; // @[RA_Mul.scala 66:39:@24.8]
  assign _GEN_3 = _T_99 ? io_A : _GEN_2; // @[RA_Mul.scala 64:39:@19.6]
  assign S_v_0 = io_eB_0[2]; // @[RA_Mul.scala 76:23:@46.4]
  assign _T_115 = io_A[15]; // @[RA_Mul.scala 77:36:@49.4]
  assign _T_116 = S_v_0 ^ _T_115; // @[RA_Mul.scala 77:30:@50.4]
  assign SC_v_0 = ~ _T_116; // @[RA_Mul.scala 77:16:@51.4]
  assign _T_119 = io_eB_1 == 3'h0; // @[RA_Mul.scala 62:19:@53.4]
  assign _T_121 = io_eB_1 == 3'h4; // @[RA_Mul.scala 62:44:@54.4]
  assign _T_122 = _T_119 | _T_121; // @[RA_Mul.scala 62:32:@55.4]
  assign _T_125 = io_eB_1 == 3'h1; // @[RA_Mul.scala 64:25:@60.6]
  assign _T_127 = io_eB_1 == 3'h2; // @[RA_Mul.scala 66:25:@65.8]
  assign _T_131 = io_eB_1 == 3'h5; // @[RA_Mul.scala 68:25:@72.10]
  assign _T_134 = io_eB_1 == 3'h6; // @[RA_Mul.scala 70:25:@78.12]
  assign _GEN_5 = _T_134 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@79.12]
  assign _GEN_6 = _T_131 ? _T_106 : _GEN_5; // @[RA_Mul.scala 68:39:@73.10]
  assign _GEN_7 = _T_127 ? _T_103 : _GEN_6; // @[RA_Mul.scala 66:39:@66.8]
  assign _GEN_8 = _T_125 ? io_A : _GEN_7; // @[RA_Mul.scala 64:39:@61.6]
  assign S_v_1 = io_eB_1[2]; // @[RA_Mul.scala 76:23:@88.4]
  assign _T_142 = S_v_1 ^ _T_115; // @[RA_Mul.scala 77:30:@92.4]
  assign SC_v_1 = ~ _T_142; // @[RA_Mul.scala 77:16:@93.4]
  assign _T_145 = io_eB_2 == 3'h0; // @[RA_Mul.scala 62:19:@95.4]
  assign _T_147 = io_eB_2 == 3'h4; // @[RA_Mul.scala 62:44:@96.4]
  assign _T_148 = _T_145 | _T_147; // @[RA_Mul.scala 62:32:@97.4]
  assign _T_151 = io_eB_2 == 3'h1; // @[RA_Mul.scala 64:25:@102.6]
  assign _T_153 = io_eB_2 == 3'h2; // @[RA_Mul.scala 66:25:@107.8]
  assign _T_157 = io_eB_2 == 3'h5; // @[RA_Mul.scala 68:25:@114.10]
  assign _T_160 = io_eB_2 == 3'h6; // @[RA_Mul.scala 70:25:@120.12]
  assign _GEN_10 = _T_160 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@121.12]
  assign _GEN_11 = _T_157 ? _T_106 : _GEN_10; // @[RA_Mul.scala 68:39:@115.10]
  assign _GEN_12 = _T_153 ? _T_103 : _GEN_11; // @[RA_Mul.scala 66:39:@108.8]
  assign _GEN_13 = _T_151 ? io_A : _GEN_12; // @[RA_Mul.scala 64:39:@103.6]
  assign S_v_2 = io_eB_2[2]; // @[RA_Mul.scala 76:23:@130.4]
  assign _T_168 = S_v_2 ^ _T_115; // @[RA_Mul.scala 77:30:@134.4]
  assign SC_v_2 = ~ _T_168; // @[RA_Mul.scala 77:16:@135.4]
  assign _T_171 = io_eB_3 == 3'h0; // @[RA_Mul.scala 62:19:@137.4]
  assign _T_173 = io_eB_3 == 3'h4; // @[RA_Mul.scala 62:44:@138.4]
  assign _T_174 = _T_171 | _T_173; // @[RA_Mul.scala 62:32:@139.4]
  assign _T_177 = io_eB_3 == 3'h1; // @[RA_Mul.scala 64:25:@144.6]
  assign _T_179 = io_eB_3 == 3'h2; // @[RA_Mul.scala 66:25:@149.8]
  assign _T_183 = io_eB_3 == 3'h5; // @[RA_Mul.scala 68:25:@156.10]
  assign _T_186 = io_eB_3 == 3'h6; // @[RA_Mul.scala 70:25:@162.12]
  assign _GEN_15 = _T_186 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@163.12]
  assign _GEN_16 = _T_183 ? _T_106 : _GEN_15; // @[RA_Mul.scala 68:39:@157.10]
  assign _GEN_17 = _T_179 ? _T_103 : _GEN_16; // @[RA_Mul.scala 66:39:@150.8]
  assign _GEN_18 = _T_177 ? io_A : _GEN_17; // @[RA_Mul.scala 64:39:@145.6]
  assign S_v_3 = io_eB_3[2]; // @[RA_Mul.scala 76:23:@172.4]
  assign _T_194 = S_v_3 ^ _T_115; // @[RA_Mul.scala 77:30:@176.4]
  assign SC_v_3 = ~ _T_194; // @[RA_Mul.scala 77:16:@177.4]
  assign _T_197 = io_eB_4 == 3'h0; // @[RA_Mul.scala 62:19:@179.4]
  assign _T_199 = io_eB_4 == 3'h4; // @[RA_Mul.scala 62:44:@180.4]
  assign _T_200 = _T_197 | _T_199; // @[RA_Mul.scala 62:32:@181.4]
  assign _T_203 = io_eB_4 == 3'h1; // @[RA_Mul.scala 64:25:@186.6]
  assign _T_205 = io_eB_4 == 3'h2; // @[RA_Mul.scala 66:25:@191.8]
  assign _T_209 = io_eB_4 == 3'h5; // @[RA_Mul.scala 68:25:@198.10]
  assign _T_212 = io_eB_4 == 3'h6; // @[RA_Mul.scala 70:25:@204.12]
  assign _GEN_20 = _T_212 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@205.12]
  assign _GEN_21 = _T_209 ? _T_106 : _GEN_20; // @[RA_Mul.scala 68:39:@199.10]
  assign _GEN_22 = _T_205 ? _T_103 : _GEN_21; // @[RA_Mul.scala 66:39:@192.8]
  assign _GEN_23 = _T_203 ? io_A : _GEN_22; // @[RA_Mul.scala 64:39:@187.6]
  assign S_v_4 = io_eB_4[2]; // @[RA_Mul.scala 76:23:@214.4]
  assign _T_220 = S_v_4 ^ _T_115; // @[RA_Mul.scala 77:30:@218.4]
  assign SC_v_4 = ~ _T_220; // @[RA_Mul.scala 77:16:@219.4]
  assign _T_223 = io_eB_5 == 3'h0; // @[RA_Mul.scala 62:19:@221.4]
  assign _T_225 = io_eB_5 == 3'h4; // @[RA_Mul.scala 62:44:@222.4]
  assign _T_226 = _T_223 | _T_225; // @[RA_Mul.scala 62:32:@223.4]
  assign _T_229 = io_eB_5 == 3'h1; // @[RA_Mul.scala 64:25:@228.6]
  assign _T_231 = io_eB_5 == 3'h2; // @[RA_Mul.scala 66:25:@233.8]
  assign _T_235 = io_eB_5 == 3'h5; // @[RA_Mul.scala 68:25:@240.10]
  assign _T_238 = io_eB_5 == 3'h6; // @[RA_Mul.scala 70:25:@246.12]
  assign _GEN_25 = _T_238 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@247.12]
  assign _GEN_26 = _T_235 ? _T_106 : _GEN_25; // @[RA_Mul.scala 68:39:@241.10]
  assign _GEN_27 = _T_231 ? _T_103 : _GEN_26; // @[RA_Mul.scala 66:39:@234.8]
  assign _GEN_28 = _T_229 ? io_A : _GEN_27; // @[RA_Mul.scala 64:39:@229.6]
  assign S_v_5 = io_eB_5[2]; // @[RA_Mul.scala 76:23:@256.4]
  assign _T_246 = S_v_5 ^ _T_115; // @[RA_Mul.scala 77:30:@260.4]
  assign SC_v_5 = ~ _T_246; // @[RA_Mul.scala 77:16:@261.4]
  assign _T_249 = io_eB_6 == 3'h0; // @[RA_Mul.scala 62:19:@263.4]
  assign _T_251 = io_eB_6 == 3'h4; // @[RA_Mul.scala 62:44:@264.4]
  assign _T_252 = _T_249 | _T_251; // @[RA_Mul.scala 62:32:@265.4]
  assign _T_255 = io_eB_6 == 3'h1; // @[RA_Mul.scala 64:25:@270.6]
  assign _T_257 = io_eB_6 == 3'h2; // @[RA_Mul.scala 66:25:@275.8]
  assign _T_261 = io_eB_6 == 3'h5; // @[RA_Mul.scala 68:25:@282.10]
  assign _T_264 = io_eB_6 == 3'h6; // @[RA_Mul.scala 70:25:@288.12]
  assign _GEN_30 = _T_264 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@289.12]
  assign _GEN_31 = _T_261 ? _T_106 : _GEN_30; // @[RA_Mul.scala 68:39:@283.10]
  assign _GEN_32 = _T_257 ? _T_103 : _GEN_31; // @[RA_Mul.scala 66:39:@276.8]
  assign _GEN_33 = _T_255 ? io_A : _GEN_32; // @[RA_Mul.scala 64:39:@271.6]
  assign S_v_6 = io_eB_6[2]; // @[RA_Mul.scala 76:23:@298.4]
  assign _T_272 = S_v_6 ^ _T_115; // @[RA_Mul.scala 77:30:@302.4]
  assign SC_v_6 = ~ _T_272; // @[RA_Mul.scala 77:16:@303.4]
  assign _T_275 = io_eB_7 == 3'h0; // @[RA_Mul.scala 62:19:@305.4]
  assign _T_277 = io_eB_7 == 3'h4; // @[RA_Mul.scala 62:44:@306.4]
  assign _T_278 = _T_275 | _T_277; // @[RA_Mul.scala 62:32:@307.4]
  assign _T_281 = io_eB_7 == 3'h1; // @[RA_Mul.scala 64:25:@312.6]
  assign _T_283 = io_eB_7 == 3'h2; // @[RA_Mul.scala 66:25:@317.8]
  assign _T_287 = io_eB_7 == 3'h5; // @[RA_Mul.scala 68:25:@324.10]
  assign _T_290 = io_eB_7 == 3'h6; // @[RA_Mul.scala 70:25:@330.12]
  assign _GEN_35 = _T_290 ? _T_111 : 16'h0; // @[RA_Mul.scala 70:38:@331.12]
  assign _GEN_36 = _T_287 ? _T_106 : _GEN_35; // @[RA_Mul.scala 68:39:@325.10]
  assign _GEN_37 = _T_283 ? _T_103 : _GEN_36; // @[RA_Mul.scala 66:39:@318.8]
  assign _GEN_38 = _T_281 ? io_A : _GEN_37; // @[RA_Mul.scala 64:39:@313.6]
  assign S_v_7 = io_eB_7[2]; // @[RA_Mul.scala 76:23:@340.4]
  assign _T_298 = S_v_7 ^ _T_115; // @[RA_Mul.scala 77:30:@344.4]
  assign SC_v_7 = ~ _T_298; // @[RA_Mul.scala 77:16:@345.4]
  assign _T_300 = {S_v_1,S_v_0}; // @[RA_Mul.scala 79:21:@347.4]
  assign _T_301 = {S_v_3,S_v_2}; // @[RA_Mul.scala 79:21:@348.4]
  assign _T_302 = {_T_301,_T_300}; // @[RA_Mul.scala 79:21:@349.4]
  assign _T_303 = {S_v_5,S_v_4}; // @[RA_Mul.scala 79:21:@350.4]
  assign _T_304 = {S_v_7,S_v_6}; // @[RA_Mul.scala 79:21:@351.4]
  assign _T_305 = {_T_304,_T_303}; // @[RA_Mul.scala 79:21:@352.4]
  assign _T_307 = {SC_v_1,SC_v_0}; // @[RA_Mul.scala 80:23:@355.4]
  assign _T_308 = {SC_v_3,SC_v_2}; // @[RA_Mul.scala 80:23:@356.4]
  assign _T_309 = {_T_308,_T_307}; // @[RA_Mul.scala 80:23:@357.4]
  assign _T_310 = {SC_v_5,SC_v_4}; // @[RA_Mul.scala 80:23:@358.4]
  assign _T_311 = {SC_v_7,SC_v_6}; // @[RA_Mul.scala 80:23:@359.4]
  assign _T_312 = {_T_311,_T_310}; // @[RA_Mul.scala 80:23:@360.4]
  assign io_PP_0 = _T_96 ? 16'h0 : _GEN_3; // @[RA_Mul.scala 63:16:@15.6 RA_Mul.scala 65:16:@20.8 RA_Mul.scala 67:16:@27.10 RA_Mul.scala 69:16:@33.12 RA_Mul.scala 71:16:@41.14 RA_Mul.scala 73:16:@44.14]
  assign io_PP_1 = _T_122 ? 16'h0 : _GEN_8; // @[RA_Mul.scala 63:16:@57.6 RA_Mul.scala 65:16:@62.8 RA_Mul.scala 67:16:@69.10 RA_Mul.scala 69:16:@75.12 RA_Mul.scala 71:16:@83.14 RA_Mul.scala 73:16:@86.14]
  assign io_PP_2 = _T_148 ? 16'h0 : _GEN_13; // @[RA_Mul.scala 63:16:@99.6 RA_Mul.scala 65:16:@104.8 RA_Mul.scala 67:16:@111.10 RA_Mul.scala 69:16:@117.12 RA_Mul.scala 71:16:@125.14 RA_Mul.scala 73:16:@128.14]
  assign io_PP_3 = _T_174 ? 16'h0 : _GEN_18; // @[RA_Mul.scala 63:16:@141.6 RA_Mul.scala 65:16:@146.8 RA_Mul.scala 67:16:@153.10 RA_Mul.scala 69:16:@159.12 RA_Mul.scala 71:16:@167.14 RA_Mul.scala 73:16:@170.14]
  assign io_PP_4 = _T_200 ? 16'h0 : _GEN_23; // @[RA_Mul.scala 63:16:@183.6 RA_Mul.scala 65:16:@188.8 RA_Mul.scala 67:16:@195.10 RA_Mul.scala 69:16:@201.12 RA_Mul.scala 71:16:@209.14 RA_Mul.scala 73:16:@212.14]
  assign io_PP_5 = _T_226 ? 16'h0 : _GEN_28; // @[RA_Mul.scala 63:16:@225.6 RA_Mul.scala 65:16:@230.8 RA_Mul.scala 67:16:@237.10 RA_Mul.scala 69:16:@243.12 RA_Mul.scala 71:16:@251.14 RA_Mul.scala 73:16:@254.14]
  assign io_PP_6 = _T_252 ? 16'h0 : _GEN_33; // @[RA_Mul.scala 63:16:@267.6 RA_Mul.scala 65:16:@272.8 RA_Mul.scala 67:16:@279.10 RA_Mul.scala 69:16:@285.12 RA_Mul.scala 71:16:@293.14 RA_Mul.scala 73:16:@296.14]
  assign io_PP_7 = _T_278 ? 16'h0 : _GEN_38; // @[RA_Mul.scala 63:16:@309.6 RA_Mul.scala 65:16:@314.8 RA_Mul.scala 67:16:@321.10 RA_Mul.scala 69:16:@327.12 RA_Mul.scala 71:16:@335.14 RA_Mul.scala 73:16:@338.14]
  assign io_SS = 8'hab; // @[RA_Mul.scala 58:9:@8.4]
  assign io_SC = {_T_312,_T_309}; // @[RA_Mul.scala 80:9:@362.4]
  assign io_S = {_T_305,_T_302}; // @[RA_Mul.scala 79:8:@354.4]
endmodule
