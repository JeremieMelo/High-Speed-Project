module BoothEncoder_radix4( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [2:0]  io_eB_0, // @[:@6.4]
  output [2:0]  io_eB_1, // @[:@6.4]
  output [2:0]  io_eB_2, // @[:@6.4]
  output [2:0]  io_eB_3, // @[:@6.4]
  output [2:0]  io_eB_4, // @[:@6.4]
  output [2:0]  io_eB_5, // @[:@6.4]
  output [2:0]  io_eB_6, // @[:@6.4]
  output [2:0]  io_eB_7, // @[:@6.4]
  input  [15:0] io_B // @[:@6.4]
);
  wire  _T_33; // @[RA_Mul.scala 36:28:@8.4]
  wire  _T_34; // @[RA_Mul.scala 36:28:@9.4]
  wire  _T_35; // @[RA_Mul.scala 36:28:@10.4]
  wire  _T_36; // @[RA_Mul.scala 36:28:@11.4]
  wire  _T_37; // @[RA_Mul.scala 36:28:@12.4]
  wire  _T_38; // @[RA_Mul.scala 36:28:@13.4]
  wire  _T_39; // @[RA_Mul.scala 36:28:@14.4]
  wire  _T_40; // @[RA_Mul.scala 36:28:@15.4]
  wire  _T_41; // @[RA_Mul.scala 36:28:@16.4]
  wire  _T_42; // @[RA_Mul.scala 36:28:@17.4]
  wire  _T_43; // @[RA_Mul.scala 36:28:@18.4]
  wire  _T_44; // @[RA_Mul.scala 36:28:@19.4]
  wire  _T_45; // @[RA_Mul.scala 36:28:@20.4]
  wire  _T_46; // @[RA_Mul.scala 36:28:@21.4]
  wire  _T_47; // @[RA_Mul.scala 36:28:@22.4]
  wire  _T_48; // @[RA_Mul.scala 36:28:@23.4]
  wire [1:0] _T_74; // @[RA_Mul.scala 36:51:@42.4]
  wire [1:0] _T_75; // @[RA_Mul.scala 36:51:@43.4]
  wire [3:0] _T_76; // @[RA_Mul.scala 36:51:@44.4]
  wire [1:0] _T_77; // @[RA_Mul.scala 36:51:@45.4]
  wire [1:0] _T_78; // @[RA_Mul.scala 36:51:@46.4]
  wire [3:0] _T_79; // @[RA_Mul.scala 36:51:@47.4]
  wire [7:0] _T_80; // @[RA_Mul.scala 36:51:@48.4]
  wire [1:0] _T_81; // @[RA_Mul.scala 36:51:@49.4]
  wire [1:0] _T_82; // @[RA_Mul.scala 36:51:@50.4]
  wire [3:0] _T_83; // @[RA_Mul.scala 36:51:@51.4]
  wire [1:0] _T_84; // @[RA_Mul.scala 36:51:@52.4]
  wire [1:0] _T_85; // @[RA_Mul.scala 36:51:@53.4]
  wire [2:0] _T_86; // @[RA_Mul.scala 36:51:@54.4]
  wire [4:0] _T_87; // @[RA_Mul.scala 36:51:@55.4]
  wire [8:0] _T_88; // @[RA_Mul.scala 36:51:@56.4]
  wire [16:0] B_ext; // @[RA_Mul.scala 36:51:@57.4]
  wire  _T_98; // @[RA_Mul.scala 41:24:@59.4]
  wire  _T_99; // @[RA_Mul.scala 41:37:@60.4]
  wire  _T_100; // @[RA_Mul.scala 41:30:@61.4]
  wire  _T_101; // @[RA_Mul.scala 42:25:@63.4]
  wire  _T_103; // @[RA_Mul.scala 42:36:@65.4]
  wire  _T_104; // @[RA_Mul.scala 42:33:@66.4]
  wire  _T_106; // @[RA_Mul.scala 42:54:@68.4]
  wire  _T_107; // @[RA_Mul.scala 42:51:@69.4]
  wire  _T_109; // @[RA_Mul.scala 42:70:@71.4]
  wire  _T_111; // @[RA_Mul.scala 42:85:@73.4]
  wire  _T_113; // @[RA_Mul.scala 42:100:@75.4]
  wire  _T_114; // @[RA_Mul.scala 42:66:@76.4]
  wire [1:0] _T_116; // @[RA_Mul.scala 44:25:@80.4]
  wire  _T_129; // @[RA_Mul.scala 41:30:@86.4]
  wire  _T_130; // @[RA_Mul.scala 42:25:@88.4]
  wire  _T_133; // @[RA_Mul.scala 42:33:@91.4]
  wire  _T_136; // @[RA_Mul.scala 42:51:@94.4]
  wire  _T_138; // @[RA_Mul.scala 42:70:@96.4]
  wire  _T_140; // @[RA_Mul.scala 42:85:@98.4]
  wire  _T_142; // @[RA_Mul.scala 42:100:@100.4]
  wire  _T_143; // @[RA_Mul.scala 42:66:@101.4]
  wire [1:0] _T_145; // @[RA_Mul.scala 44:25:@105.4]
  wire  _T_158; // @[RA_Mul.scala 41:30:@111.4]
  wire  _T_159; // @[RA_Mul.scala 42:25:@113.4]
  wire  _T_162; // @[RA_Mul.scala 42:33:@116.4]
  wire  _T_165; // @[RA_Mul.scala 42:51:@119.4]
  wire  _T_167; // @[RA_Mul.scala 42:70:@121.4]
  wire  _T_169; // @[RA_Mul.scala 42:85:@123.4]
  wire  _T_171; // @[RA_Mul.scala 42:100:@125.4]
  wire  _T_172; // @[RA_Mul.scala 42:66:@126.4]
  wire [1:0] _T_174; // @[RA_Mul.scala 44:25:@130.4]
  wire  _T_187; // @[RA_Mul.scala 41:30:@136.4]
  wire  _T_188; // @[RA_Mul.scala 42:25:@138.4]
  wire  _T_191; // @[RA_Mul.scala 42:33:@141.4]
  wire  _T_194; // @[RA_Mul.scala 42:51:@144.4]
  wire  _T_196; // @[RA_Mul.scala 42:70:@146.4]
  wire  _T_198; // @[RA_Mul.scala 42:85:@148.4]
  wire  _T_200; // @[RA_Mul.scala 42:100:@150.4]
  wire  _T_201; // @[RA_Mul.scala 42:66:@151.4]
  wire [1:0] _T_203; // @[RA_Mul.scala 44:25:@155.4]
  wire  _T_216; // @[RA_Mul.scala 41:30:@161.4]
  wire  _T_217; // @[RA_Mul.scala 42:25:@163.4]
  wire  _T_220; // @[RA_Mul.scala 42:33:@166.4]
  wire  _T_223; // @[RA_Mul.scala 42:51:@169.4]
  wire  _T_225; // @[RA_Mul.scala 42:70:@171.4]
  wire  _T_227; // @[RA_Mul.scala 42:85:@173.4]
  wire  _T_229; // @[RA_Mul.scala 42:100:@175.4]
  wire  _T_230; // @[RA_Mul.scala 42:66:@176.4]
  wire [1:0] _T_232; // @[RA_Mul.scala 44:25:@180.4]
  wire  _T_245; // @[RA_Mul.scala 41:30:@186.4]
  wire  _T_246; // @[RA_Mul.scala 42:25:@188.4]
  wire  _T_249; // @[RA_Mul.scala 42:33:@191.4]
  wire  _T_252; // @[RA_Mul.scala 42:51:@194.4]
  wire  _T_254; // @[RA_Mul.scala 42:70:@196.4]
  wire  _T_256; // @[RA_Mul.scala 42:85:@198.4]
  wire  _T_258; // @[RA_Mul.scala 42:100:@200.4]
  wire  _T_259; // @[RA_Mul.scala 42:66:@201.4]
  wire [1:0] _T_261; // @[RA_Mul.scala 44:25:@205.4]
  wire  _T_274; // @[RA_Mul.scala 41:30:@211.4]
  wire  _T_275; // @[RA_Mul.scala 42:25:@213.4]
  wire  _T_278; // @[RA_Mul.scala 42:33:@216.4]
  wire  _T_281; // @[RA_Mul.scala 42:51:@219.4]
  wire  _T_283; // @[RA_Mul.scala 42:70:@221.4]
  wire  _T_285; // @[RA_Mul.scala 42:85:@223.4]
  wire  _T_287; // @[RA_Mul.scala 42:100:@225.4]
  wire  _T_288; // @[RA_Mul.scala 42:66:@226.4]
  wire [1:0] _T_290; // @[RA_Mul.scala 44:25:@230.4]
  wire  _T_303; // @[RA_Mul.scala 41:30:@236.4]
  wire  _T_304; // @[RA_Mul.scala 42:25:@238.4]
  wire  _T_307; // @[RA_Mul.scala 42:33:@241.4]
  wire  _T_310; // @[RA_Mul.scala 42:51:@244.4]
  wire  _T_312; // @[RA_Mul.scala 42:70:@246.4]
  wire  _T_314; // @[RA_Mul.scala 42:85:@248.4]
  wire  _T_316; // @[RA_Mul.scala 42:100:@250.4]
  wire  _T_317; // @[RA_Mul.scala 42:66:@251.4]
  wire [1:0] _T_319; // @[RA_Mul.scala 44:25:@255.4]
  assign _T_33 = io_B[0]; // @[RA_Mul.scala 36:28:@8.4]
  assign _T_34 = io_B[1]; // @[RA_Mul.scala 36:28:@9.4]
  assign _T_35 = io_B[2]; // @[RA_Mul.scala 36:28:@10.4]
  assign _T_36 = io_B[3]; // @[RA_Mul.scala 36:28:@11.4]
  assign _T_37 = io_B[4]; // @[RA_Mul.scala 36:28:@12.4]
  assign _T_38 = io_B[5]; // @[RA_Mul.scala 36:28:@13.4]
  assign _T_39 = io_B[6]; // @[RA_Mul.scala 36:28:@14.4]
  assign _T_40 = io_B[7]; // @[RA_Mul.scala 36:28:@15.4]
  assign _T_41 = io_B[8]; // @[RA_Mul.scala 36:28:@16.4]
  assign _T_42 = io_B[9]; // @[RA_Mul.scala 36:28:@17.4]
  assign _T_43 = io_B[10]; // @[RA_Mul.scala 36:28:@18.4]
  assign _T_44 = io_B[11]; // @[RA_Mul.scala 36:28:@19.4]
  assign _T_45 = io_B[12]; // @[RA_Mul.scala 36:28:@20.4]
  assign _T_46 = io_B[13]; // @[RA_Mul.scala 36:28:@21.4]
  assign _T_47 = io_B[14]; // @[RA_Mul.scala 36:28:@22.4]
  assign _T_48 = io_B[15]; // @[RA_Mul.scala 36:28:@23.4]
  assign _T_74 = {_T_34,_T_33}; // @[RA_Mul.scala 36:51:@42.4]
  assign _T_75 = {_T_36,_T_35}; // @[RA_Mul.scala 36:51:@43.4]
  assign _T_76 = {_T_75,_T_74}; // @[RA_Mul.scala 36:51:@44.4]
  assign _T_77 = {_T_38,_T_37}; // @[RA_Mul.scala 36:51:@45.4]
  assign _T_78 = {_T_40,_T_39}; // @[RA_Mul.scala 36:51:@46.4]
  assign _T_79 = {_T_78,_T_77}; // @[RA_Mul.scala 36:51:@47.4]
  assign _T_80 = {_T_79,_T_76}; // @[RA_Mul.scala 36:51:@48.4]
  assign _T_81 = {_T_42,_T_41}; // @[RA_Mul.scala 36:51:@49.4]
  assign _T_82 = {_T_44,_T_43}; // @[RA_Mul.scala 36:51:@50.4]
  assign _T_83 = {_T_82,_T_81}; // @[RA_Mul.scala 36:51:@51.4]
  assign _T_84 = {_T_46,_T_45}; // @[RA_Mul.scala 36:51:@52.4]
  assign _T_85 = {1'h0,_T_48}; // @[RA_Mul.scala 36:51:@53.4]
  assign _T_86 = {_T_85,_T_47}; // @[RA_Mul.scala 36:51:@54.4]
  assign _T_87 = {_T_86,_T_84}; // @[RA_Mul.scala 36:51:@55.4]
  assign _T_88 = {_T_87,_T_83}; // @[RA_Mul.scala 36:51:@56.4]
  assign B_ext = {_T_88,_T_80}; // @[RA_Mul.scala 36:51:@57.4]
  assign _T_98 = B_ext[1]; // @[RA_Mul.scala 41:24:@59.4]
  assign _T_99 = B_ext[0]; // @[RA_Mul.scala 41:37:@60.4]
  assign _T_100 = _T_98 ^ _T_99; // @[RA_Mul.scala 41:30:@61.4]
  assign _T_101 = B_ext[2]; // @[RA_Mul.scala 42:25:@63.4]
  assign _T_103 = ~ _T_98; // @[RA_Mul.scala 42:36:@65.4]
  assign _T_104 = _T_101 & _T_103; // @[RA_Mul.scala 42:33:@66.4]
  assign _T_106 = ~ _T_99; // @[RA_Mul.scala 42:54:@68.4]
  assign _T_107 = _T_104 & _T_106; // @[RA_Mul.scala 42:51:@69.4]
  assign _T_109 = ~ _T_101; // @[RA_Mul.scala 42:70:@71.4]
  assign _T_111 = _T_109 & _T_98; // @[RA_Mul.scala 42:85:@73.4]
  assign _T_113 = _T_111 & _T_99; // @[RA_Mul.scala 42:100:@75.4]
  assign _T_114 = _T_107 | _T_113; // @[RA_Mul.scala 42:66:@76.4]
  assign _T_116 = {_T_101,_T_114}; // @[RA_Mul.scala 44:25:@80.4]
  assign _T_129 = _T_101 ^ _T_98; // @[RA_Mul.scala 41:30:@86.4]
  assign _T_130 = B_ext[3]; // @[RA_Mul.scala 42:25:@88.4]
  assign _T_133 = _T_130 & _T_109; // @[RA_Mul.scala 42:33:@91.4]
  assign _T_136 = _T_133 & _T_103; // @[RA_Mul.scala 42:51:@94.4]
  assign _T_138 = ~ _T_130; // @[RA_Mul.scala 42:70:@96.4]
  assign _T_140 = _T_138 & _T_101; // @[RA_Mul.scala 42:85:@98.4]
  assign _T_142 = _T_140 & _T_98; // @[RA_Mul.scala 42:100:@100.4]
  assign _T_143 = _T_136 | _T_142; // @[RA_Mul.scala 42:66:@101.4]
  assign _T_145 = {_T_130,_T_143}; // @[RA_Mul.scala 44:25:@105.4]
  assign _T_158 = _T_130 ^ _T_101; // @[RA_Mul.scala 41:30:@111.4]
  assign _T_159 = B_ext[4]; // @[RA_Mul.scala 42:25:@113.4]
  assign _T_162 = _T_159 & _T_138; // @[RA_Mul.scala 42:33:@116.4]
  assign _T_165 = _T_162 & _T_109; // @[RA_Mul.scala 42:51:@119.4]
  assign _T_167 = ~ _T_159; // @[RA_Mul.scala 42:70:@121.4]
  assign _T_169 = _T_167 & _T_130; // @[RA_Mul.scala 42:85:@123.4]
  assign _T_171 = _T_169 & _T_101; // @[RA_Mul.scala 42:100:@125.4]
  assign _T_172 = _T_165 | _T_171; // @[RA_Mul.scala 42:66:@126.4]
  assign _T_174 = {_T_159,_T_172}; // @[RA_Mul.scala 44:25:@130.4]
  assign _T_187 = _T_159 ^ _T_130; // @[RA_Mul.scala 41:30:@136.4]
  assign _T_188 = B_ext[5]; // @[RA_Mul.scala 42:25:@138.4]
  assign _T_191 = _T_188 & _T_167; // @[RA_Mul.scala 42:33:@141.4]
  assign _T_194 = _T_191 & _T_138; // @[RA_Mul.scala 42:51:@144.4]
  assign _T_196 = ~ _T_188; // @[RA_Mul.scala 42:70:@146.4]
  assign _T_198 = _T_196 & _T_159; // @[RA_Mul.scala 42:85:@148.4]
  assign _T_200 = _T_198 & _T_130; // @[RA_Mul.scala 42:100:@150.4]
  assign _T_201 = _T_194 | _T_200; // @[RA_Mul.scala 42:66:@151.4]
  assign _T_203 = {_T_188,_T_201}; // @[RA_Mul.scala 44:25:@155.4]
  assign _T_216 = _T_188 ^ _T_159; // @[RA_Mul.scala 41:30:@161.4]
  assign _T_217 = B_ext[6]; // @[RA_Mul.scala 42:25:@163.4]
  assign _T_220 = _T_217 & _T_196; // @[RA_Mul.scala 42:33:@166.4]
  assign _T_223 = _T_220 & _T_167; // @[RA_Mul.scala 42:51:@169.4]
  assign _T_225 = ~ _T_217; // @[RA_Mul.scala 42:70:@171.4]
  assign _T_227 = _T_225 & _T_188; // @[RA_Mul.scala 42:85:@173.4]
  assign _T_229 = _T_227 & _T_159; // @[RA_Mul.scala 42:100:@175.4]
  assign _T_230 = _T_223 | _T_229; // @[RA_Mul.scala 42:66:@176.4]
  assign _T_232 = {_T_217,_T_230}; // @[RA_Mul.scala 44:25:@180.4]
  assign _T_245 = _T_217 ^ _T_188; // @[RA_Mul.scala 41:30:@186.4]
  assign _T_246 = B_ext[7]; // @[RA_Mul.scala 42:25:@188.4]
  assign _T_249 = _T_246 & _T_225; // @[RA_Mul.scala 42:33:@191.4]
  assign _T_252 = _T_249 & _T_196; // @[RA_Mul.scala 42:51:@194.4]
  assign _T_254 = ~ _T_246; // @[RA_Mul.scala 42:70:@196.4]
  assign _T_256 = _T_254 & _T_217; // @[RA_Mul.scala 42:85:@198.4]
  assign _T_258 = _T_256 & _T_188; // @[RA_Mul.scala 42:100:@200.4]
  assign _T_259 = _T_252 | _T_258; // @[RA_Mul.scala 42:66:@201.4]
  assign _T_261 = {_T_246,_T_259}; // @[RA_Mul.scala 44:25:@205.4]
  assign _T_274 = _T_246 ^ _T_217; // @[RA_Mul.scala 41:30:@211.4]
  assign _T_275 = B_ext[8]; // @[RA_Mul.scala 42:25:@213.4]
  assign _T_278 = _T_275 & _T_254; // @[RA_Mul.scala 42:33:@216.4]
  assign _T_281 = _T_278 & _T_225; // @[RA_Mul.scala 42:51:@219.4]
  assign _T_283 = ~ _T_275; // @[RA_Mul.scala 42:70:@221.4]
  assign _T_285 = _T_283 & _T_246; // @[RA_Mul.scala 42:85:@223.4]
  assign _T_287 = _T_285 & _T_217; // @[RA_Mul.scala 42:100:@225.4]
  assign _T_288 = _T_281 | _T_287; // @[RA_Mul.scala 42:66:@226.4]
  assign _T_290 = {_T_275,_T_288}; // @[RA_Mul.scala 44:25:@230.4]
  assign _T_303 = _T_275 ^ _T_246; // @[RA_Mul.scala 41:30:@236.4]
  assign _T_304 = B_ext[9]; // @[RA_Mul.scala 42:25:@238.4]
  assign _T_307 = _T_304 & _T_283; // @[RA_Mul.scala 42:33:@241.4]
  assign _T_310 = _T_307 & _T_254; // @[RA_Mul.scala 42:51:@244.4]
  assign _T_312 = ~ _T_304; // @[RA_Mul.scala 42:70:@246.4]
  assign _T_314 = _T_312 & _T_275; // @[RA_Mul.scala 42:85:@248.4]
  assign _T_316 = _T_314 & _T_246; // @[RA_Mul.scala 42:100:@250.4]
  assign _T_317 = _T_310 | _T_316; // @[RA_Mul.scala 42:66:@251.4]
  assign _T_319 = {_T_304,_T_317}; // @[RA_Mul.scala 44:25:@255.4]
  assign io_eB_0 = {_T_116,_T_100}; // @[RA_Mul.scala 44:15:@82.4]
  assign io_eB_1 = {_T_145,_T_129}; // @[RA_Mul.scala 44:15:@107.4]
  assign io_eB_2 = {_T_174,_T_158}; // @[RA_Mul.scala 44:15:@132.4]
  assign io_eB_3 = {_T_203,_T_187}; // @[RA_Mul.scala 44:15:@157.4]
  assign io_eB_4 = {_T_232,_T_216}; // @[RA_Mul.scala 44:15:@182.4]
  assign io_eB_5 = {_T_261,_T_245}; // @[RA_Mul.scala 44:15:@207.4]
  assign io_eB_6 = {_T_290,_T_274}; // @[RA_Mul.scala 44:15:@232.4]
  assign io_eB_7 = {_T_319,_T_303}; // @[RA_Mul.scala 44:15:@257.4]
endmodule
