module HA( // @[:@3.2]
  output  io_s, // @[:@6.4]
  output  io_cout, // @[:@6.4]
  input   io_a, // @[:@6.4]
  input   io_b // @[:@6.4]
);
  assign io_s = io_a ^ io_b; // @[RA_Mul.scala 12:8:@11.4]
  assign io_cout = io_a & io_b; // @[RA_Mul.scala 11:11:@9.4]
endmodule
module FA( // @[:@13.2]
  output  io_s, // @[:@16.4]
  output  io_cout, // @[:@16.4]
  input   io_a, // @[:@16.4]
  input   io_b, // @[:@16.4]
  input   io_cin // @[:@16.4]
);
  wire  _T_15; // @[RA_Mul.scala 35:16:@18.4]
  wire  _T_17; // @[RA_Mul.scala 36:20:@21.4]
  wire  _T_18; // @[RA_Mul.scala 36:36:@22.4]
  wire  _T_19; // @[RA_Mul.scala 36:28:@23.4]
  wire  _T_20; // @[RA_Mul.scala 36:54:@24.4]
  assign _T_15 = io_a ^ io_b; // @[RA_Mul.scala 35:16:@18.4]
  assign _T_17 = io_a & io_b; // @[RA_Mul.scala 36:20:@21.4]
  assign _T_18 = io_a & io_cin; // @[RA_Mul.scala 36:36:@22.4]
  assign _T_19 = _T_17 | _T_18; // @[RA_Mul.scala 36:28:@23.4]
  assign _T_20 = io_b & io_cin; // @[RA_Mul.scala 36:54:@24.4]
  assign io_s = _T_15 ^ io_cin; // @[RA_Mul.scala 35:8:@20.4]
  assign io_cout = _T_19 | _T_20; // @[RA_Mul.scala 36:11:@26.4]
endmodule
module Reduction_2( // @[:@478.2]
  input   clock, // @[:@479.4]
  input   reset, // @[:@480.4]
  output  io_matrix_o_0_0, // @[:@481.4]
  output  io_matrix_o_0_1, // @[:@481.4]
  output  io_matrix_o_0_2, // @[:@481.4]
  output  io_matrix_o_0_3, // @[:@481.4]
  output  io_matrix_o_0_4, // @[:@481.4]
  output  io_matrix_o_0_5, // @[:@481.4]
  output  io_matrix_o_0_6, // @[:@481.4]
  output  io_matrix_o_0_7, // @[:@481.4]
  output  io_matrix_o_0_8, // @[:@481.4]
  output  io_matrix_o_0_9, // @[:@481.4]
  output  io_matrix_o_0_10, // @[:@481.4]
  output  io_matrix_o_0_11, // @[:@481.4]
  output  io_matrix_o_0_12, // @[:@481.4]
  output  io_matrix_o_0_13, // @[:@481.4]
  output  io_matrix_o_0_14, // @[:@481.4]
  output  io_matrix_o_0_15, // @[:@481.4]
  output  io_matrix_o_0_16, // @[:@481.4]
  output  io_matrix_o_0_17, // @[:@481.4]
  output  io_matrix_o_0_18, // @[:@481.4]
  output  io_matrix_o_0_19, // @[:@481.4]
  output  io_matrix_o_0_20, // @[:@481.4]
  output  io_matrix_o_0_21, // @[:@481.4]
  output  io_matrix_o_0_22, // @[:@481.4]
  output  io_matrix_o_0_23, // @[:@481.4]
  output  io_matrix_o_0_24, // @[:@481.4]
  output  io_matrix_o_0_25, // @[:@481.4]
  output  io_matrix_o_0_26, // @[:@481.4]
  output  io_matrix_o_0_27, // @[:@481.4]
  output  io_matrix_o_0_28, // @[:@481.4]
  output  io_matrix_o_0_29, // @[:@481.4]
  output  io_matrix_o_0_30, // @[:@481.4]
  output  io_matrix_o_0_31, // @[:@481.4]
  output  io_matrix_o_1_0, // @[:@481.4]
  output  io_matrix_o_1_1, // @[:@481.4]
  output  io_matrix_o_1_2, // @[:@481.4]
  output  io_matrix_o_1_3, // @[:@481.4]
  output  io_matrix_o_1_4, // @[:@481.4]
  output  io_matrix_o_1_5, // @[:@481.4]
  output  io_matrix_o_1_6, // @[:@481.4]
  output  io_matrix_o_1_7, // @[:@481.4]
  output  io_matrix_o_1_8, // @[:@481.4]
  output  io_matrix_o_1_9, // @[:@481.4]
  output  io_matrix_o_1_10, // @[:@481.4]
  output  io_matrix_o_1_11, // @[:@481.4]
  output  io_matrix_o_1_12, // @[:@481.4]
  output  io_matrix_o_1_13, // @[:@481.4]
  output  io_matrix_o_1_14, // @[:@481.4]
  output  io_matrix_o_1_15, // @[:@481.4]
  output  io_matrix_o_1_16, // @[:@481.4]
  output  io_matrix_o_1_17, // @[:@481.4]
  output  io_matrix_o_1_18, // @[:@481.4]
  output  io_matrix_o_1_19, // @[:@481.4]
  output  io_matrix_o_1_20, // @[:@481.4]
  output  io_matrix_o_1_21, // @[:@481.4]
  output  io_matrix_o_1_22, // @[:@481.4]
  output  io_matrix_o_1_23, // @[:@481.4]
  output  io_matrix_o_1_24, // @[:@481.4]
  output  io_matrix_o_1_25, // @[:@481.4]
  output  io_matrix_o_1_26, // @[:@481.4]
  output  io_matrix_o_1_27, // @[:@481.4]
  output  io_matrix_o_1_28, // @[:@481.4]
  output  io_matrix_o_1_29, // @[:@481.4]
  output  io_matrix_o_1_30, // @[:@481.4]
  output  io_matrix_o_1_31, // @[:@481.4]
  output  io_matrix_o_2_0, // @[:@481.4]
  output  io_matrix_o_2_1, // @[:@481.4]
  output  io_matrix_o_2_2, // @[:@481.4]
  output  io_matrix_o_2_3, // @[:@481.4]
  output  io_matrix_o_2_4, // @[:@481.4]
  output  io_matrix_o_2_5, // @[:@481.4]
  output  io_matrix_o_2_6, // @[:@481.4]
  output  io_matrix_o_2_7, // @[:@481.4]
  output  io_matrix_o_2_8, // @[:@481.4]
  output  io_matrix_o_2_9, // @[:@481.4]
  output  io_matrix_o_2_10, // @[:@481.4]
  output  io_matrix_o_2_11, // @[:@481.4]
  output  io_matrix_o_2_12, // @[:@481.4]
  output  io_matrix_o_2_13, // @[:@481.4]
  output  io_matrix_o_2_14, // @[:@481.4]
  output  io_matrix_o_2_15, // @[:@481.4]
  output  io_matrix_o_2_16, // @[:@481.4]
  output  io_matrix_o_2_17, // @[:@481.4]
  output  io_matrix_o_2_18, // @[:@481.4]
  output  io_matrix_o_2_19, // @[:@481.4]
  output  io_matrix_o_2_20, // @[:@481.4]
  output  io_matrix_o_2_21, // @[:@481.4]
  output  io_matrix_o_2_22, // @[:@481.4]
  output  io_matrix_o_2_23, // @[:@481.4]
  output  io_matrix_o_2_24, // @[:@481.4]
  output  io_matrix_o_2_25, // @[:@481.4]
  output  io_matrix_o_2_26, // @[:@481.4]
  output  io_matrix_o_2_27, // @[:@481.4]
  output  io_matrix_o_2_28, // @[:@481.4]
  output  io_matrix_o_2_29, // @[:@481.4]
  output  io_matrix_o_2_30, // @[:@481.4]
  output  io_matrix_o_2_31, // @[:@481.4]
  output  io_matrix_o_3_0, // @[:@481.4]
  output  io_matrix_o_3_1, // @[:@481.4]
  output  io_matrix_o_3_2, // @[:@481.4]
  output  io_matrix_o_3_3, // @[:@481.4]
  output  io_matrix_o_3_4, // @[:@481.4]
  output  io_matrix_o_3_5, // @[:@481.4]
  output  io_matrix_o_3_6, // @[:@481.4]
  output  io_matrix_o_3_7, // @[:@481.4]
  output  io_matrix_o_3_8, // @[:@481.4]
  output  io_matrix_o_3_9, // @[:@481.4]
  output  io_matrix_o_3_10, // @[:@481.4]
  output  io_matrix_o_3_11, // @[:@481.4]
  output  io_matrix_o_3_12, // @[:@481.4]
  output  io_matrix_o_3_13, // @[:@481.4]
  output  io_matrix_o_3_14, // @[:@481.4]
  output  io_matrix_o_3_15, // @[:@481.4]
  output  io_matrix_o_3_16, // @[:@481.4]
  output  io_matrix_o_3_17, // @[:@481.4]
  output  io_matrix_o_3_18, // @[:@481.4]
  output  io_matrix_o_3_19, // @[:@481.4]
  output  io_matrix_o_3_20, // @[:@481.4]
  output  io_matrix_o_3_21, // @[:@481.4]
  output  io_matrix_o_3_22, // @[:@481.4]
  output  io_matrix_o_3_23, // @[:@481.4]
  output  io_matrix_o_3_24, // @[:@481.4]
  output  io_matrix_o_3_25, // @[:@481.4]
  output  io_matrix_o_3_26, // @[:@481.4]
  output  io_matrix_o_3_27, // @[:@481.4]
  output  io_matrix_o_3_28, // @[:@481.4]
  output  io_matrix_o_3_29, // @[:@481.4]
  output  io_matrix_o_3_30, // @[:@481.4]
  output  io_matrix_o_3_31, // @[:@481.4]
  input   io_matrix_i_0_0, // @[:@481.4]
  input   io_matrix_i_0_1, // @[:@481.4]
  input   io_matrix_i_0_2, // @[:@481.4]
  input   io_matrix_i_0_3, // @[:@481.4]
  input   io_matrix_i_0_4, // @[:@481.4]
  input   io_matrix_i_0_5, // @[:@481.4]
  input   io_matrix_i_0_6, // @[:@481.4]
  input   io_matrix_i_0_7, // @[:@481.4]
  input   io_matrix_i_0_8, // @[:@481.4]
  input   io_matrix_i_0_9, // @[:@481.4]
  input   io_matrix_i_0_10, // @[:@481.4]
  input   io_matrix_i_0_11, // @[:@481.4]
  input   io_matrix_i_0_12, // @[:@481.4]
  input   io_matrix_i_0_13, // @[:@481.4]
  input   io_matrix_i_0_14, // @[:@481.4]
  input   io_matrix_i_0_15, // @[:@481.4]
  input   io_matrix_i_0_16, // @[:@481.4]
  input   io_matrix_i_0_17, // @[:@481.4]
  input   io_matrix_i_0_18, // @[:@481.4]
  input   io_matrix_i_0_19, // @[:@481.4]
  input   io_matrix_i_0_20, // @[:@481.4]
  input   io_matrix_i_0_21, // @[:@481.4]
  input   io_matrix_i_0_22, // @[:@481.4]
  input   io_matrix_i_0_23, // @[:@481.4]
  input   io_matrix_i_0_24, // @[:@481.4]
  input   io_matrix_i_0_25, // @[:@481.4]
  input   io_matrix_i_0_26, // @[:@481.4]
  input   io_matrix_i_0_27, // @[:@481.4]
  input   io_matrix_i_0_28, // @[:@481.4]
  input   io_matrix_i_0_29, // @[:@481.4]
  input   io_matrix_i_0_30, // @[:@481.4]
  input   io_matrix_i_0_31, // @[:@481.4]
  input   io_matrix_i_1_0, // @[:@481.4]
  input   io_matrix_i_1_1, // @[:@481.4]
  input   io_matrix_i_1_2, // @[:@481.4]
  input   io_matrix_i_1_3, // @[:@481.4]
  input   io_matrix_i_1_4, // @[:@481.4]
  input   io_matrix_i_1_5, // @[:@481.4]
  input   io_matrix_i_1_6, // @[:@481.4]
  input   io_matrix_i_1_7, // @[:@481.4]
  input   io_matrix_i_1_8, // @[:@481.4]
  input   io_matrix_i_1_9, // @[:@481.4]
  input   io_matrix_i_1_10, // @[:@481.4]
  input   io_matrix_i_1_11, // @[:@481.4]
  input   io_matrix_i_1_12, // @[:@481.4]
  input   io_matrix_i_1_13, // @[:@481.4]
  input   io_matrix_i_1_14, // @[:@481.4]
  input   io_matrix_i_1_15, // @[:@481.4]
  input   io_matrix_i_1_16, // @[:@481.4]
  input   io_matrix_i_1_17, // @[:@481.4]
  input   io_matrix_i_1_18, // @[:@481.4]
  input   io_matrix_i_1_19, // @[:@481.4]
  input   io_matrix_i_1_20, // @[:@481.4]
  input   io_matrix_i_1_21, // @[:@481.4]
  input   io_matrix_i_1_22, // @[:@481.4]
  input   io_matrix_i_1_23, // @[:@481.4]
  input   io_matrix_i_1_24, // @[:@481.4]
  input   io_matrix_i_1_25, // @[:@481.4]
  input   io_matrix_i_1_26, // @[:@481.4]
  input   io_matrix_i_1_27, // @[:@481.4]
  input   io_matrix_i_1_28, // @[:@481.4]
  input   io_matrix_i_1_29, // @[:@481.4]
  input   io_matrix_i_1_30, // @[:@481.4]
  input   io_matrix_i_1_31, // @[:@481.4]
  input   io_matrix_i_2_0, // @[:@481.4]
  input   io_matrix_i_2_1, // @[:@481.4]
  input   io_matrix_i_2_2, // @[:@481.4]
  input   io_matrix_i_2_3, // @[:@481.4]
  input   io_matrix_i_2_4, // @[:@481.4]
  input   io_matrix_i_2_5, // @[:@481.4]
  input   io_matrix_i_2_6, // @[:@481.4]
  input   io_matrix_i_2_7, // @[:@481.4]
  input   io_matrix_i_2_8, // @[:@481.4]
  input   io_matrix_i_2_9, // @[:@481.4]
  input   io_matrix_i_2_10, // @[:@481.4]
  input   io_matrix_i_2_11, // @[:@481.4]
  input   io_matrix_i_2_12, // @[:@481.4]
  input   io_matrix_i_2_13, // @[:@481.4]
  input   io_matrix_i_2_14, // @[:@481.4]
  input   io_matrix_i_2_15, // @[:@481.4]
  input   io_matrix_i_2_16, // @[:@481.4]
  input   io_matrix_i_2_17, // @[:@481.4]
  input   io_matrix_i_2_18, // @[:@481.4]
  input   io_matrix_i_2_19, // @[:@481.4]
  input   io_matrix_i_2_20, // @[:@481.4]
  input   io_matrix_i_2_21, // @[:@481.4]
  input   io_matrix_i_2_22, // @[:@481.4]
  input   io_matrix_i_2_23, // @[:@481.4]
  input   io_matrix_i_2_24, // @[:@481.4]
  input   io_matrix_i_2_25, // @[:@481.4]
  input   io_matrix_i_2_26, // @[:@481.4]
  input   io_matrix_i_2_27, // @[:@481.4]
  input   io_matrix_i_2_28, // @[:@481.4]
  input   io_matrix_i_2_29, // @[:@481.4]
  input   io_matrix_i_2_30, // @[:@481.4]
  input   io_matrix_i_2_31, // @[:@481.4]
  input   io_matrix_i_3_0, // @[:@481.4]
  input   io_matrix_i_3_1, // @[:@481.4]
  input   io_matrix_i_3_2, // @[:@481.4]
  input   io_matrix_i_3_3, // @[:@481.4]
  input   io_matrix_i_3_4, // @[:@481.4]
  input   io_matrix_i_3_5, // @[:@481.4]
  input   io_matrix_i_3_6, // @[:@481.4]
  input   io_matrix_i_3_7, // @[:@481.4]
  input   io_matrix_i_3_8, // @[:@481.4]
  input   io_matrix_i_3_9, // @[:@481.4]
  input   io_matrix_i_3_10, // @[:@481.4]
  input   io_matrix_i_3_11, // @[:@481.4]
  input   io_matrix_i_3_12, // @[:@481.4]
  input   io_matrix_i_3_13, // @[:@481.4]
  input   io_matrix_i_3_14, // @[:@481.4]
  input   io_matrix_i_3_15, // @[:@481.4]
  input   io_matrix_i_3_16, // @[:@481.4]
  input   io_matrix_i_3_17, // @[:@481.4]
  input   io_matrix_i_3_18, // @[:@481.4]
  input   io_matrix_i_3_19, // @[:@481.4]
  input   io_matrix_i_3_20, // @[:@481.4]
  input   io_matrix_i_3_21, // @[:@481.4]
  input   io_matrix_i_3_22, // @[:@481.4]
  input   io_matrix_i_3_23, // @[:@481.4]
  input   io_matrix_i_3_24, // @[:@481.4]
  input   io_matrix_i_3_25, // @[:@481.4]
  input   io_matrix_i_3_26, // @[:@481.4]
  input   io_matrix_i_3_27, // @[:@481.4]
  input   io_matrix_i_3_28, // @[:@481.4]
  input   io_matrix_i_3_29, // @[:@481.4]
  input   io_matrix_i_3_30, // @[:@481.4]
  input   io_matrix_i_3_31, // @[:@481.4]
  input   io_matrix_i_4_0, // @[:@481.4]
  input   io_matrix_i_4_1, // @[:@481.4]
  input   io_matrix_i_4_2, // @[:@481.4]
  input   io_matrix_i_4_3, // @[:@481.4]
  input   io_matrix_i_4_4, // @[:@481.4]
  input   io_matrix_i_4_5, // @[:@481.4]
  input   io_matrix_i_4_6, // @[:@481.4]
  input   io_matrix_i_4_7, // @[:@481.4]
  input   io_matrix_i_4_8, // @[:@481.4]
  input   io_matrix_i_4_9, // @[:@481.4]
  input   io_matrix_i_4_10, // @[:@481.4]
  input   io_matrix_i_4_11, // @[:@481.4]
  input   io_matrix_i_4_12, // @[:@481.4]
  input   io_matrix_i_4_13, // @[:@481.4]
  input   io_matrix_i_4_14, // @[:@481.4]
  input   io_matrix_i_4_15, // @[:@481.4]
  input   io_matrix_i_4_16, // @[:@481.4]
  input   io_matrix_i_4_17, // @[:@481.4]
  input   io_matrix_i_4_18, // @[:@481.4]
  input   io_matrix_i_4_19, // @[:@481.4]
  input   io_matrix_i_4_20, // @[:@481.4]
  input   io_matrix_i_4_21, // @[:@481.4]
  input   io_matrix_i_4_22, // @[:@481.4]
  input   io_matrix_i_4_23, // @[:@481.4]
  input   io_matrix_i_4_24, // @[:@481.4]
  input   io_matrix_i_4_25, // @[:@481.4]
  input   io_matrix_i_4_26, // @[:@481.4]
  input   io_matrix_i_4_27, // @[:@481.4]
  input   io_matrix_i_4_28, // @[:@481.4]
  input   io_matrix_i_4_29, // @[:@481.4]
  input   io_matrix_i_4_30, // @[:@481.4]
  input   io_matrix_i_4_31, // @[:@481.4]
  input   io_matrix_i_5_0, // @[:@481.4]
  input   io_matrix_i_5_1, // @[:@481.4]
  input   io_matrix_i_5_2, // @[:@481.4]
  input   io_matrix_i_5_3, // @[:@481.4]
  input   io_matrix_i_5_4, // @[:@481.4]
  input   io_matrix_i_5_5, // @[:@481.4]
  input   io_matrix_i_5_6, // @[:@481.4]
  input   io_matrix_i_5_7, // @[:@481.4]
  input   io_matrix_i_5_8, // @[:@481.4]
  input   io_matrix_i_5_9, // @[:@481.4]
  input   io_matrix_i_5_10, // @[:@481.4]
  input   io_matrix_i_5_11, // @[:@481.4]
  input   io_matrix_i_5_12, // @[:@481.4]
  input   io_matrix_i_5_13, // @[:@481.4]
  input   io_matrix_i_5_14, // @[:@481.4]
  input   io_matrix_i_5_15, // @[:@481.4]
  input   io_matrix_i_5_16, // @[:@481.4]
  input   io_matrix_i_5_17, // @[:@481.4]
  input   io_matrix_i_5_18, // @[:@481.4]
  input   io_matrix_i_5_19, // @[:@481.4]
  input   io_matrix_i_5_20, // @[:@481.4]
  input   io_matrix_i_5_21, // @[:@481.4]
  input   io_matrix_i_5_22, // @[:@481.4]
  input   io_matrix_i_5_23, // @[:@481.4]
  input   io_matrix_i_5_24, // @[:@481.4]
  input   io_matrix_i_5_25, // @[:@481.4]
  input   io_matrix_i_5_26, // @[:@481.4]
  input   io_matrix_i_5_27, // @[:@481.4]
  input   io_matrix_i_5_28, // @[:@481.4]
  input   io_matrix_i_5_29, // @[:@481.4]
  input   io_matrix_i_5_30, // @[:@481.4]
  input   io_matrix_i_5_31 // @[:@481.4]
);
  wire  HA_io_s; // @[RA_Mul.scala 18:21:@487.4]
  wire  HA_io_cout; // @[RA_Mul.scala 18:21:@487.4]
  wire  HA_io_a; // @[RA_Mul.scala 18:21:@487.4]
  wire  HA_io_b; // @[RA_Mul.scala 18:21:@487.4]
  wire  FA_io_s; // @[RA_Mul.scala 42:21:@501.4]
  wire  FA_io_cout; // @[RA_Mul.scala 42:21:@501.4]
  wire  FA_io_a; // @[RA_Mul.scala 42:21:@501.4]
  wire  FA_io_b; // @[RA_Mul.scala 42:21:@501.4]
  wire  FA_io_cin; // @[RA_Mul.scala 42:21:@501.4]
  wire  FA_1_io_s; // @[RA_Mul.scala 42:21:@520.4]
  wire  FA_1_io_cout; // @[RA_Mul.scala 42:21:@520.4]
  wire  FA_1_io_a; // @[RA_Mul.scala 42:21:@520.4]
  wire  FA_1_io_b; // @[RA_Mul.scala 42:21:@520.4]
  wire  FA_1_io_cin; // @[RA_Mul.scala 42:21:@520.4]
  wire  FA_2_io_s; // @[RA_Mul.scala 42:21:@531.4]
  wire  FA_2_io_cout; // @[RA_Mul.scala 42:21:@531.4]
  wire  FA_2_io_a; // @[RA_Mul.scala 42:21:@531.4]
  wire  FA_2_io_b; // @[RA_Mul.scala 42:21:@531.4]
  wire  FA_2_io_cin; // @[RA_Mul.scala 42:21:@531.4]
  wire  FA_3_io_s; // @[RA_Mul.scala 42:21:@541.4]
  wire  FA_3_io_cout; // @[RA_Mul.scala 42:21:@541.4]
  wire  FA_3_io_a; // @[RA_Mul.scala 42:21:@541.4]
  wire  FA_3_io_b; // @[RA_Mul.scala 42:21:@541.4]
  wire  FA_3_io_cin; // @[RA_Mul.scala 42:21:@541.4]
  wire  FA_4_io_s; // @[RA_Mul.scala 42:21:@551.4]
  wire  FA_4_io_cout; // @[RA_Mul.scala 42:21:@551.4]
  wire  FA_4_io_a; // @[RA_Mul.scala 42:21:@551.4]
  wire  FA_4_io_b; // @[RA_Mul.scala 42:21:@551.4]
  wire  FA_4_io_cin; // @[RA_Mul.scala 42:21:@551.4]
  wire  FA_5_io_s; // @[RA_Mul.scala 42:21:@561.4]
  wire  FA_5_io_cout; // @[RA_Mul.scala 42:21:@561.4]
  wire  FA_5_io_a; // @[RA_Mul.scala 42:21:@561.4]
  wire  FA_5_io_b; // @[RA_Mul.scala 42:21:@561.4]
  wire  FA_5_io_cin; // @[RA_Mul.scala 42:21:@561.4]
  wire  FA_6_io_s; // @[RA_Mul.scala 42:21:@571.4]
  wire  FA_6_io_cout; // @[RA_Mul.scala 42:21:@571.4]
  wire  FA_6_io_a; // @[RA_Mul.scala 42:21:@571.4]
  wire  FA_6_io_b; // @[RA_Mul.scala 42:21:@571.4]
  wire  FA_6_io_cin; // @[RA_Mul.scala 42:21:@571.4]
  wire  FA_7_io_s; // @[RA_Mul.scala 42:21:@581.4]
  wire  FA_7_io_cout; // @[RA_Mul.scala 42:21:@581.4]
  wire  FA_7_io_a; // @[RA_Mul.scala 42:21:@581.4]
  wire  FA_7_io_b; // @[RA_Mul.scala 42:21:@581.4]
  wire  FA_7_io_cin; // @[RA_Mul.scala 42:21:@581.4]
  wire  FA_8_io_s; // @[RA_Mul.scala 42:21:@589.4]
  wire  FA_8_io_cout; // @[RA_Mul.scala 42:21:@589.4]
  wire  FA_8_io_a; // @[RA_Mul.scala 42:21:@589.4]
  wire  FA_8_io_b; // @[RA_Mul.scala 42:21:@589.4]
  wire  FA_8_io_cin; // @[RA_Mul.scala 42:21:@589.4]
  wire  FA_9_io_s; // @[RA_Mul.scala 42:21:@598.4]
  wire  FA_9_io_cout; // @[RA_Mul.scala 42:21:@598.4]
  wire  FA_9_io_a; // @[RA_Mul.scala 42:21:@598.4]
  wire  FA_9_io_b; // @[RA_Mul.scala 42:21:@598.4]
  wire  FA_9_io_cin; // @[RA_Mul.scala 42:21:@598.4]
  wire  HA_1_io_s; // @[RA_Mul.scala 18:21:@606.4]
  wire  HA_1_io_cout; // @[RA_Mul.scala 18:21:@606.4]
  wire  HA_1_io_a; // @[RA_Mul.scala 18:21:@606.4]
  wire  HA_1_io_b; // @[RA_Mul.scala 18:21:@606.4]
  wire  FA_10_io_s; // @[RA_Mul.scala 42:21:@613.4]
  wire  FA_10_io_cout; // @[RA_Mul.scala 42:21:@613.4]
  wire  FA_10_io_a; // @[RA_Mul.scala 42:21:@613.4]
  wire  FA_10_io_b; // @[RA_Mul.scala 42:21:@613.4]
  wire  FA_10_io_cin; // @[RA_Mul.scala 42:21:@613.4]
  wire  HA_2_io_s; // @[RA_Mul.scala 18:21:@621.4]
  wire  HA_2_io_cout; // @[RA_Mul.scala 18:21:@621.4]
  wire  HA_2_io_a; // @[RA_Mul.scala 18:21:@621.4]
  wire  HA_2_io_b; // @[RA_Mul.scala 18:21:@621.4]
  wire  FA_11_io_s; // @[RA_Mul.scala 42:21:@628.4]
  wire  FA_11_io_cout; // @[RA_Mul.scala 42:21:@628.4]
  wire  FA_11_io_a; // @[RA_Mul.scala 42:21:@628.4]
  wire  FA_11_io_b; // @[RA_Mul.scala 42:21:@628.4]
  wire  FA_11_io_cin; // @[RA_Mul.scala 42:21:@628.4]
  wire  FA_12_io_s; // @[RA_Mul.scala 42:21:@636.4]
  wire  FA_12_io_cout; // @[RA_Mul.scala 42:21:@636.4]
  wire  FA_12_io_a; // @[RA_Mul.scala 42:21:@636.4]
  wire  FA_12_io_b; // @[RA_Mul.scala 42:21:@636.4]
  wire  FA_12_io_cin; // @[RA_Mul.scala 42:21:@636.4]
  wire  FA_13_io_s; // @[RA_Mul.scala 42:21:@644.4]
  wire  FA_13_io_cout; // @[RA_Mul.scala 42:21:@644.4]
  wire  FA_13_io_a; // @[RA_Mul.scala 42:21:@644.4]
  wire  FA_13_io_b; // @[RA_Mul.scala 42:21:@644.4]
  wire  FA_13_io_cin; // @[RA_Mul.scala 42:21:@644.4]
  wire  FA_14_io_s; // @[RA_Mul.scala 42:21:@652.4]
  wire  FA_14_io_cout; // @[RA_Mul.scala 42:21:@652.4]
  wire  FA_14_io_a; // @[RA_Mul.scala 42:21:@652.4]
  wire  FA_14_io_b; // @[RA_Mul.scala 42:21:@652.4]
  wire  FA_14_io_cin; // @[RA_Mul.scala 42:21:@652.4]
  wire  FA_15_io_s; // @[RA_Mul.scala 42:21:@660.4]
  wire  FA_15_io_cout; // @[RA_Mul.scala 42:21:@660.4]
  wire  FA_15_io_a; // @[RA_Mul.scala 42:21:@660.4]
  wire  FA_15_io_b; // @[RA_Mul.scala 42:21:@660.4]
  wire  FA_15_io_cin; // @[RA_Mul.scala 42:21:@660.4]
  wire  FA_16_io_s; // @[RA_Mul.scala 42:21:@668.4]
  wire  FA_16_io_cout; // @[RA_Mul.scala 42:21:@668.4]
  wire  FA_16_io_a; // @[RA_Mul.scala 42:21:@668.4]
  wire  FA_16_io_b; // @[RA_Mul.scala 42:21:@668.4]
  wire  FA_16_io_cin; // @[RA_Mul.scala 42:21:@668.4]
  wire  FA_17_io_s; // @[RA_Mul.scala 42:21:@676.4]
  wire  FA_17_io_cout; // @[RA_Mul.scala 42:21:@676.4]
  wire  FA_17_io_a; // @[RA_Mul.scala 42:21:@676.4]
  wire  FA_17_io_b; // @[RA_Mul.scala 42:21:@676.4]
  wire  FA_17_io_cin; // @[RA_Mul.scala 42:21:@676.4]
  wire  FA_18_io_s; // @[RA_Mul.scala 42:21:@684.4]
  wire  FA_18_io_cout; // @[RA_Mul.scala 42:21:@684.4]
  wire  FA_18_io_a; // @[RA_Mul.scala 42:21:@684.4]
  wire  FA_18_io_b; // @[RA_Mul.scala 42:21:@684.4]
  wire  FA_18_io_cin; // @[RA_Mul.scala 42:21:@684.4]
  wire  FA_19_io_s; // @[RA_Mul.scala 42:21:@692.4]
  wire  FA_19_io_cout; // @[RA_Mul.scala 42:21:@692.4]
  wire  FA_19_io_a; // @[RA_Mul.scala 42:21:@692.4]
  wire  FA_19_io_b; // @[RA_Mul.scala 42:21:@692.4]
  wire  FA_19_io_cin; // @[RA_Mul.scala 42:21:@692.4]
  wire  FA_20_io_s; // @[RA_Mul.scala 42:21:@700.4]
  wire  FA_20_io_cout; // @[RA_Mul.scala 42:21:@700.4]
  wire  FA_20_io_a; // @[RA_Mul.scala 42:21:@700.4]
  wire  FA_20_io_b; // @[RA_Mul.scala 42:21:@700.4]
  wire  FA_20_io_cin; // @[RA_Mul.scala 42:21:@700.4]
  wire  FA_21_io_s; // @[RA_Mul.scala 42:21:@708.4]
  wire  FA_21_io_cout; // @[RA_Mul.scala 42:21:@708.4]
  wire  FA_21_io_a; // @[RA_Mul.scala 42:21:@708.4]
  wire  FA_21_io_b; // @[RA_Mul.scala 42:21:@708.4]
  wire  FA_21_io_cin; // @[RA_Mul.scala 42:21:@708.4]
  wire  HA_3_io_s; // @[RA_Mul.scala 18:21:@716.4]
  wire  HA_3_io_cout; // @[RA_Mul.scala 18:21:@716.4]
  wire  HA_3_io_a; // @[RA_Mul.scala 18:21:@716.4]
  wire  HA_3_io_b; // @[RA_Mul.scala 18:21:@716.4]
  wire  FA_22_io_s; // @[RA_Mul.scala 42:21:@723.4]
  wire  FA_22_io_cout; // @[RA_Mul.scala 42:21:@723.4]
  wire  FA_22_io_a; // @[RA_Mul.scala 42:21:@723.4]
  wire  FA_22_io_b; // @[RA_Mul.scala 42:21:@723.4]
  wire  FA_22_io_cin; // @[RA_Mul.scala 42:21:@723.4]
  wire  FA_23_io_s; // @[RA_Mul.scala 42:21:@732.4]
  wire  FA_23_io_cout; // @[RA_Mul.scala 42:21:@732.4]
  wire  FA_23_io_a; // @[RA_Mul.scala 42:21:@732.4]
  wire  FA_23_io_b; // @[RA_Mul.scala 42:21:@732.4]
  wire  FA_23_io_cin; // @[RA_Mul.scala 42:21:@732.4]
  wire  FA_24_io_s; // @[RA_Mul.scala 42:21:@742.4]
  wire  FA_24_io_cout; // @[RA_Mul.scala 42:21:@742.4]
  wire  FA_24_io_a; // @[RA_Mul.scala 42:21:@742.4]
  wire  FA_24_io_b; // @[RA_Mul.scala 42:21:@742.4]
  wire  FA_24_io_cin; // @[RA_Mul.scala 42:21:@742.4]
  wire  FA_25_io_s; // @[RA_Mul.scala 42:21:@752.4]
  wire  FA_25_io_cout; // @[RA_Mul.scala 42:21:@752.4]
  wire  FA_25_io_a; // @[RA_Mul.scala 42:21:@752.4]
  wire  FA_25_io_b; // @[RA_Mul.scala 42:21:@752.4]
  wire  FA_25_io_cin; // @[RA_Mul.scala 42:21:@752.4]
  wire  FA_26_io_s; // @[RA_Mul.scala 42:21:@762.4]
  wire  FA_26_io_cout; // @[RA_Mul.scala 42:21:@762.4]
  wire  FA_26_io_a; // @[RA_Mul.scala 42:21:@762.4]
  wire  FA_26_io_b; // @[RA_Mul.scala 42:21:@762.4]
  wire  FA_26_io_cin; // @[RA_Mul.scala 42:21:@762.4]
  wire  FA_27_io_s; // @[RA_Mul.scala 42:21:@772.4]
  wire  FA_27_io_cout; // @[RA_Mul.scala 42:21:@772.4]
  wire  FA_27_io_a; // @[RA_Mul.scala 42:21:@772.4]
  wire  FA_27_io_b; // @[RA_Mul.scala 42:21:@772.4]
  wire  FA_27_io_cin; // @[RA_Mul.scala 42:21:@772.4]
  wire  FA_28_io_s; // @[RA_Mul.scala 42:21:@789.4]
  wire  FA_28_io_cout; // @[RA_Mul.scala 42:21:@789.4]
  wire  FA_28_io_a; // @[RA_Mul.scala 42:21:@789.4]
  wire  FA_28_io_b; // @[RA_Mul.scala 42:21:@789.4]
  wire  FA_28_io_cin; // @[RA_Mul.scala 42:21:@789.4]
  HA HA ( // @[RA_Mul.scala 18:21:@487.4]
    .io_s(HA_io_s),
    .io_cout(HA_io_cout),
    .io_a(HA_io_a),
    .io_b(HA_io_b)
  );
  FA FA ( // @[RA_Mul.scala 42:21:@501.4]
    .io_s(FA_io_s),
    .io_cout(FA_io_cout),
    .io_a(FA_io_a),
    .io_b(FA_io_b),
    .io_cin(FA_io_cin)
  );
  FA FA_1 ( // @[RA_Mul.scala 42:21:@520.4]
    .io_s(FA_1_io_s),
    .io_cout(FA_1_io_cout),
    .io_a(FA_1_io_a),
    .io_b(FA_1_io_b),
    .io_cin(FA_1_io_cin)
  );
  FA FA_2 ( // @[RA_Mul.scala 42:21:@531.4]
    .io_s(FA_2_io_s),
    .io_cout(FA_2_io_cout),
    .io_a(FA_2_io_a),
    .io_b(FA_2_io_b),
    .io_cin(FA_2_io_cin)
  );
  FA FA_3 ( // @[RA_Mul.scala 42:21:@541.4]
    .io_s(FA_3_io_s),
    .io_cout(FA_3_io_cout),
    .io_a(FA_3_io_a),
    .io_b(FA_3_io_b),
    .io_cin(FA_3_io_cin)
  );
  FA FA_4 ( // @[RA_Mul.scala 42:21:@551.4]
    .io_s(FA_4_io_s),
    .io_cout(FA_4_io_cout),
    .io_a(FA_4_io_a),
    .io_b(FA_4_io_b),
    .io_cin(FA_4_io_cin)
  );
  FA FA_5 ( // @[RA_Mul.scala 42:21:@561.4]
    .io_s(FA_5_io_s),
    .io_cout(FA_5_io_cout),
    .io_a(FA_5_io_a),
    .io_b(FA_5_io_b),
    .io_cin(FA_5_io_cin)
  );
  FA FA_6 ( // @[RA_Mul.scala 42:21:@571.4]
    .io_s(FA_6_io_s),
    .io_cout(FA_6_io_cout),
    .io_a(FA_6_io_a),
    .io_b(FA_6_io_b),
    .io_cin(FA_6_io_cin)
  );
  FA FA_7 ( // @[RA_Mul.scala 42:21:@581.4]
    .io_s(FA_7_io_s),
    .io_cout(FA_7_io_cout),
    .io_a(FA_7_io_a),
    .io_b(FA_7_io_b),
    .io_cin(FA_7_io_cin)
  );
  FA FA_8 ( // @[RA_Mul.scala 42:21:@589.4]
    .io_s(FA_8_io_s),
    .io_cout(FA_8_io_cout),
    .io_a(FA_8_io_a),
    .io_b(FA_8_io_b),
    .io_cin(FA_8_io_cin)
  );
  FA FA_9 ( // @[RA_Mul.scala 42:21:@598.4]
    .io_s(FA_9_io_s),
    .io_cout(FA_9_io_cout),
    .io_a(FA_9_io_a),
    .io_b(FA_9_io_b),
    .io_cin(FA_9_io_cin)
  );
  HA HA_1 ( // @[RA_Mul.scala 18:21:@606.4]
    .io_s(HA_1_io_s),
    .io_cout(HA_1_io_cout),
    .io_a(HA_1_io_a),
    .io_b(HA_1_io_b)
  );
  FA FA_10 ( // @[RA_Mul.scala 42:21:@613.4]
    .io_s(FA_10_io_s),
    .io_cout(FA_10_io_cout),
    .io_a(FA_10_io_a),
    .io_b(FA_10_io_b),
    .io_cin(FA_10_io_cin)
  );
  HA HA_2 ( // @[RA_Mul.scala 18:21:@621.4]
    .io_s(HA_2_io_s),
    .io_cout(HA_2_io_cout),
    .io_a(HA_2_io_a),
    .io_b(HA_2_io_b)
  );
  FA FA_11 ( // @[RA_Mul.scala 42:21:@628.4]
    .io_s(FA_11_io_s),
    .io_cout(FA_11_io_cout),
    .io_a(FA_11_io_a),
    .io_b(FA_11_io_b),
    .io_cin(FA_11_io_cin)
  );
  FA FA_12 ( // @[RA_Mul.scala 42:21:@636.4]
    .io_s(FA_12_io_s),
    .io_cout(FA_12_io_cout),
    .io_a(FA_12_io_a),
    .io_b(FA_12_io_b),
    .io_cin(FA_12_io_cin)
  );
  FA FA_13 ( // @[RA_Mul.scala 42:21:@644.4]
    .io_s(FA_13_io_s),
    .io_cout(FA_13_io_cout),
    .io_a(FA_13_io_a),
    .io_b(FA_13_io_b),
    .io_cin(FA_13_io_cin)
  );
  FA FA_14 ( // @[RA_Mul.scala 42:21:@652.4]
    .io_s(FA_14_io_s),
    .io_cout(FA_14_io_cout),
    .io_a(FA_14_io_a),
    .io_b(FA_14_io_b),
    .io_cin(FA_14_io_cin)
  );
  FA FA_15 ( // @[RA_Mul.scala 42:21:@660.4]
    .io_s(FA_15_io_s),
    .io_cout(FA_15_io_cout),
    .io_a(FA_15_io_a),
    .io_b(FA_15_io_b),
    .io_cin(FA_15_io_cin)
  );
  FA FA_16 ( // @[RA_Mul.scala 42:21:@668.4]
    .io_s(FA_16_io_s),
    .io_cout(FA_16_io_cout),
    .io_a(FA_16_io_a),
    .io_b(FA_16_io_b),
    .io_cin(FA_16_io_cin)
  );
  FA FA_17 ( // @[RA_Mul.scala 42:21:@676.4]
    .io_s(FA_17_io_s),
    .io_cout(FA_17_io_cout),
    .io_a(FA_17_io_a),
    .io_b(FA_17_io_b),
    .io_cin(FA_17_io_cin)
  );
  FA FA_18 ( // @[RA_Mul.scala 42:21:@684.4]
    .io_s(FA_18_io_s),
    .io_cout(FA_18_io_cout),
    .io_a(FA_18_io_a),
    .io_b(FA_18_io_b),
    .io_cin(FA_18_io_cin)
  );
  FA FA_19 ( // @[RA_Mul.scala 42:21:@692.4]
    .io_s(FA_19_io_s),
    .io_cout(FA_19_io_cout),
    .io_a(FA_19_io_a),
    .io_b(FA_19_io_b),
    .io_cin(FA_19_io_cin)
  );
  FA FA_20 ( // @[RA_Mul.scala 42:21:@700.4]
    .io_s(FA_20_io_s),
    .io_cout(FA_20_io_cout),
    .io_a(FA_20_io_a),
    .io_b(FA_20_io_b),
    .io_cin(FA_20_io_cin)
  );
  FA FA_21 ( // @[RA_Mul.scala 42:21:@708.4]
    .io_s(FA_21_io_s),
    .io_cout(FA_21_io_cout),
    .io_a(FA_21_io_a),
    .io_b(FA_21_io_b),
    .io_cin(FA_21_io_cin)
  );
  HA HA_3 ( // @[RA_Mul.scala 18:21:@716.4]
    .io_s(HA_3_io_s),
    .io_cout(HA_3_io_cout),
    .io_a(HA_3_io_a),
    .io_b(HA_3_io_b)
  );
  FA FA_22 ( // @[RA_Mul.scala 42:21:@723.4]
    .io_s(FA_22_io_s),
    .io_cout(FA_22_io_cout),
    .io_a(FA_22_io_a),
    .io_b(FA_22_io_b),
    .io_cin(FA_22_io_cin)
  );
  FA FA_23 ( // @[RA_Mul.scala 42:21:@732.4]
    .io_s(FA_23_io_s),
    .io_cout(FA_23_io_cout),
    .io_a(FA_23_io_a),
    .io_b(FA_23_io_b),
    .io_cin(FA_23_io_cin)
  );
  FA FA_24 ( // @[RA_Mul.scala 42:21:@742.4]
    .io_s(FA_24_io_s),
    .io_cout(FA_24_io_cout),
    .io_a(FA_24_io_a),
    .io_b(FA_24_io_b),
    .io_cin(FA_24_io_cin)
  );
  FA FA_25 ( // @[RA_Mul.scala 42:21:@752.4]
    .io_s(FA_25_io_s),
    .io_cout(FA_25_io_cout),
    .io_a(FA_25_io_a),
    .io_b(FA_25_io_b),
    .io_cin(FA_25_io_cin)
  );
  FA FA_26 ( // @[RA_Mul.scala 42:21:@762.4]
    .io_s(FA_26_io_s),
    .io_cout(FA_26_io_cout),
    .io_a(FA_26_io_a),
    .io_b(FA_26_io_b),
    .io_cin(FA_26_io_cin)
  );
  FA FA_27 ( // @[RA_Mul.scala 42:21:@772.4]
    .io_s(FA_27_io_s),
    .io_cout(FA_27_io_cout),
    .io_a(FA_27_io_a),
    .io_b(FA_27_io_b),
    .io_cin(FA_27_io_cin)
  );
  FA FA_28 ( // @[RA_Mul.scala 42:21:@789.4]
    .io_s(FA_28_io_s),
    .io_cout(FA_28_io_cout),
    .io_a(FA_28_io_a),
    .io_b(FA_28_io_b),
    .io_cin(FA_28_io_cin)
  );
  assign io_matrix_o_0_0 = io_matrix_i_0_0; // @[RA_Mul.scala 297:21:@483.4]
  assign io_matrix_o_0_1 = HA_io_s; // @[RA_Mul.scala 21:7:@492.4]
  assign io_matrix_o_0_2 = io_matrix_i_0_2; // @[RA_Mul.scala 303:21:@497.4]
  assign io_matrix_o_0_3 = FA_io_s; // @[RA_Mul.scala 46:7:@507.4]
  assign io_matrix_o_0_4 = io_matrix_i_0_4; // @[RA_Mul.scala 309:21:@512.4]
  assign io_matrix_o_0_5 = io_matrix_i_0_5; // @[RA_Mul.scala 313:21:@516.4]
  assign io_matrix_o_0_6 = FA_1_io_s; // @[RA_Mul.scala 46:7:@526.4]
  assign io_matrix_o_0_7 = FA_2_io_s; // @[RA_Mul.scala 46:7:@537.4]
  assign io_matrix_o_0_8 = FA_3_io_s; // @[RA_Mul.scala 46:7:@547.4]
  assign io_matrix_o_0_9 = FA_4_io_s; // @[RA_Mul.scala 46:7:@557.4]
  assign io_matrix_o_0_10 = FA_5_io_s; // @[RA_Mul.scala 46:7:@567.4]
  assign io_matrix_o_0_11 = FA_6_io_s; // @[RA_Mul.scala 46:7:@577.4]
  assign io_matrix_o_0_12 = FA_7_io_s; // @[RA_Mul.scala 46:7:@587.4]
  assign io_matrix_o_0_13 = FA_9_io_s; // @[RA_Mul.scala 46:7:@604.4]
  assign io_matrix_o_0_14 = FA_10_io_s; // @[RA_Mul.scala 46:7:@619.4]
  assign io_matrix_o_0_15 = FA_11_io_s; // @[RA_Mul.scala 46:7:@634.4]
  assign io_matrix_o_0_16 = FA_13_io_s; // @[RA_Mul.scala 46:7:@650.4]
  assign io_matrix_o_0_17 = FA_15_io_s; // @[RA_Mul.scala 46:7:@666.4]
  assign io_matrix_o_0_18 = FA_17_io_s; // @[RA_Mul.scala 46:7:@682.4]
  assign io_matrix_o_0_19 = FA_19_io_s; // @[RA_Mul.scala 46:7:@698.4]
  assign io_matrix_o_0_20 = FA_21_io_s; // @[RA_Mul.scala 46:7:@714.4]
  assign io_matrix_o_0_21 = FA_22_io_s; // @[RA_Mul.scala 46:7:@729.4]
  assign io_matrix_o_0_22 = FA_23_io_s; // @[RA_Mul.scala 46:7:@738.4]
  assign io_matrix_o_0_23 = FA_24_io_s; // @[RA_Mul.scala 46:7:@748.4]
  assign io_matrix_o_0_24 = FA_25_io_s; // @[RA_Mul.scala 46:7:@758.4]
  assign io_matrix_o_0_25 = FA_26_io_s; // @[RA_Mul.scala 46:7:@768.4]
  assign io_matrix_o_0_26 = FA_27_io_s; // @[RA_Mul.scala 46:7:@778.4]
  assign io_matrix_o_0_27 = io_matrix_i_0_27; // @[RA_Mul.scala 378:22:@782.4]
  assign io_matrix_o_0_28 = io_matrix_i_0_28; // @[RA_Mul.scala 382:22:@785.4]
  assign io_matrix_o_0_29 = FA_28_io_s; // @[RA_Mul.scala 46:7:@795.4]
  assign io_matrix_o_0_30 = io_matrix_i_0_30; // @[RA_Mul.scala 389:22:@800.4]
  assign io_matrix_o_0_31 = io_matrix_i_0_31; // @[RA_Mul.scala 393:22:@803.4]
  assign io_matrix_o_1_0 = 1'h0; // @[RA_Mul.scala 293:19:@484.4]
  assign io_matrix_o_1_1 = 1'h0; // @[RA_Mul.scala 293:19:@494.4]
  assign io_matrix_o_1_2 = 1'h0; // @[RA_Mul.scala 22:10:@493.4 RA_Mul.scala 293:19:@498.4]
  assign io_matrix_o_1_3 = 1'h0; // @[RA_Mul.scala 293:19:@509.4]
  assign io_matrix_o_1_4 = io_matrix_i_1_4; // @[RA_Mul.scala 47:10:@508.4 RA_Mul.scala 310:21:@513.4]
  assign io_matrix_o_1_5 = io_matrix_i_1_5; // @[RA_Mul.scala 314:21:@517.4]
  assign io_matrix_o_1_6 = io_matrix_i_3_6; // @[RA_Mul.scala 318:21:@528.4]
  assign io_matrix_o_1_7 = FA_1_io_cout; // @[RA_Mul.scala 47:10:@527.4]
  assign io_matrix_o_1_8 = FA_2_io_cout; // @[RA_Mul.scala 47:10:@538.4]
  assign io_matrix_o_1_9 = FA_3_io_cout; // @[RA_Mul.scala 47:10:@548.4]
  assign io_matrix_o_1_10 = FA_4_io_cout; // @[RA_Mul.scala 47:10:@558.4]
  assign io_matrix_o_1_11 = FA_5_io_cout; // @[RA_Mul.scala 47:10:@568.4]
  assign io_matrix_o_1_12 = FA_6_io_cout; // @[RA_Mul.scala 47:10:@578.4]
  assign io_matrix_o_1_13 = FA_7_io_cout; // @[RA_Mul.scala 47:10:@588.4]
  assign io_matrix_o_1_14 = FA_9_io_cout; // @[RA_Mul.scala 47:10:@605.4]
  assign io_matrix_o_1_15 = FA_10_io_cout; // @[RA_Mul.scala 47:10:@620.4]
  assign io_matrix_o_1_16 = FA_11_io_cout; // @[RA_Mul.scala 47:10:@635.4]
  assign io_matrix_o_1_17 = FA_13_io_cout; // @[RA_Mul.scala 47:10:@651.4]
  assign io_matrix_o_1_18 = FA_15_io_cout; // @[RA_Mul.scala 47:10:@667.4]
  assign io_matrix_o_1_19 = FA_17_io_cout; // @[RA_Mul.scala 47:10:@683.4]
  assign io_matrix_o_1_20 = FA_19_io_cout; // @[RA_Mul.scala 47:10:@699.4]
  assign io_matrix_o_1_21 = FA_21_io_cout; // @[RA_Mul.scala 47:10:@715.4]
  assign io_matrix_o_1_22 = FA_22_io_cout; // @[RA_Mul.scala 47:10:@730.4]
  assign io_matrix_o_1_23 = FA_23_io_cout; // @[RA_Mul.scala 47:10:@739.4]
  assign io_matrix_o_1_24 = FA_24_io_cout; // @[RA_Mul.scala 47:10:@749.4]
  assign io_matrix_o_1_25 = FA_25_io_cout; // @[RA_Mul.scala 47:10:@759.4]
  assign io_matrix_o_1_26 = FA_26_io_cout; // @[RA_Mul.scala 47:10:@769.4]
  assign io_matrix_o_1_27 = FA_27_io_cout; // @[RA_Mul.scala 47:10:@779.4]
  assign io_matrix_o_1_28 = io_matrix_i_1_28; // @[RA_Mul.scala 383:22:@786.4]
  assign io_matrix_o_1_29 = 1'h0; // @[RA_Mul.scala 293:19:@797.4]
  assign io_matrix_o_1_30 = FA_28_io_cout; // @[RA_Mul.scala 47:10:@796.4]
  assign io_matrix_o_1_31 = 1'h0; // @[RA_Mul.scala 293:19:@804.4]
  assign io_matrix_o_2_0 = 1'h0; // @[RA_Mul.scala 293:19:@485.4]
  assign io_matrix_o_2_1 = 1'h0; // @[RA_Mul.scala 293:19:@495.4]
  assign io_matrix_o_2_2 = 1'h0; // @[RA_Mul.scala 293:19:@499.4]
  assign io_matrix_o_2_3 = 1'h0; // @[RA_Mul.scala 293:19:@510.4]
  assign io_matrix_o_2_4 = 1'h0; // @[RA_Mul.scala 293:19:@514.4]
  assign io_matrix_o_2_5 = 1'h0; // @[RA_Mul.scala 293:19:@518.4]
  assign io_matrix_o_2_6 = 1'h0; // @[RA_Mul.scala 293:19:@529.4]
  assign io_matrix_o_2_7 = 1'h0; // @[RA_Mul.scala 293:19:@539.4]
  assign io_matrix_o_2_8 = 1'h0; // @[RA_Mul.scala 293:19:@549.4]
  assign io_matrix_o_2_9 = io_matrix_i_3_9; // @[RA_Mul.scala 328:21:@559.4]
  assign io_matrix_o_2_10 = io_matrix_i_3_10; // @[RA_Mul.scala 332:22:@569.4]
  assign io_matrix_o_2_11 = io_matrix_i_3_11; // @[RA_Mul.scala 336:22:@579.4]
  assign io_matrix_o_2_12 = FA_8_io_s; // @[RA_Mul.scala 46:7:@595.4]
  assign io_matrix_o_2_13 = HA_1_io_s; // @[RA_Mul.scala 21:7:@611.4]
  assign io_matrix_o_2_14 = HA_2_io_s; // @[RA_Mul.scala 21:7:@626.4]
  assign io_matrix_o_2_15 = FA_12_io_s; // @[RA_Mul.scala 46:7:@642.4]
  assign io_matrix_o_2_16 = FA_14_io_s; // @[RA_Mul.scala 46:7:@658.4]
  assign io_matrix_o_2_17 = FA_16_io_s; // @[RA_Mul.scala 46:7:@674.4]
  assign io_matrix_o_2_18 = FA_18_io_s; // @[RA_Mul.scala 46:7:@690.4]
  assign io_matrix_o_2_19 = FA_20_io_s; // @[RA_Mul.scala 46:7:@706.4]
  assign io_matrix_o_2_20 = HA_3_io_s; // @[RA_Mul.scala 21:7:@721.4]
  assign io_matrix_o_2_21 = io_matrix_i_3_21; // @[RA_Mul.scala 358:22:@731.4]
  assign io_matrix_o_2_22 = io_matrix_i_3_22; // @[RA_Mul.scala 361:22:@740.4]
  assign io_matrix_o_2_23 = io_matrix_i_3_23; // @[RA_Mul.scala 365:22:@750.4]
  assign io_matrix_o_2_24 = io_matrix_i_3_24; // @[RA_Mul.scala 369:22:@760.4]
  assign io_matrix_o_2_25 = 1'h0; // @[RA_Mul.scala 293:19:@770.4]
  assign io_matrix_o_2_26 = 1'h0; // @[RA_Mul.scala 293:19:@780.4]
  assign io_matrix_o_2_27 = io_matrix_i_1_27; // @[RA_Mul.scala 379:22:@783.4]
  assign io_matrix_o_2_28 = 1'h0; // @[RA_Mul.scala 293:19:@787.4]
  assign io_matrix_o_2_29 = 1'h0; // @[RA_Mul.scala 293:19:@798.4]
  assign io_matrix_o_2_30 = io_matrix_i_1_30; // @[RA_Mul.scala 390:22:@801.4]
  assign io_matrix_o_2_31 = 1'h0; // @[RA_Mul.scala 293:19:@805.4]
  assign io_matrix_o_3_0 = 1'h0; // @[RA_Mul.scala 293:19:@486.4]
  assign io_matrix_o_3_1 = 1'h0; // @[RA_Mul.scala 293:19:@496.4]
  assign io_matrix_o_3_2 = 1'h0; // @[RA_Mul.scala 293:19:@500.4]
  assign io_matrix_o_3_3 = 1'h0; // @[RA_Mul.scala 293:19:@511.4]
  assign io_matrix_o_3_4 = 1'h0; // @[RA_Mul.scala 293:19:@515.4]
  assign io_matrix_o_3_5 = 1'h0; // @[RA_Mul.scala 293:19:@519.4]
  assign io_matrix_o_3_6 = 1'h0; // @[RA_Mul.scala 293:19:@530.4]
  assign io_matrix_o_3_7 = 1'h0; // @[RA_Mul.scala 293:19:@540.4]
  assign io_matrix_o_3_8 = 1'h0; // @[RA_Mul.scala 293:19:@550.4]
  assign io_matrix_o_3_9 = io_matrix_i_4_9; // @[RA_Mul.scala 329:21:@560.4]
  assign io_matrix_o_3_10 = 1'h0; // @[RA_Mul.scala 293:19:@570.4]
  assign io_matrix_o_3_11 = 1'h0; // @[RA_Mul.scala 293:19:@580.4]
  assign io_matrix_o_3_12 = 1'h0; // @[RA_Mul.scala 293:19:@597.4]
  assign io_matrix_o_3_13 = FA_8_io_cout; // @[RA_Mul.scala 47:10:@596.4]
  assign io_matrix_o_3_14 = HA_1_io_cout; // @[RA_Mul.scala 22:10:@612.4]
  assign io_matrix_o_3_15 = HA_2_io_cout; // @[RA_Mul.scala 22:10:@627.4]
  assign io_matrix_o_3_16 = FA_12_io_cout; // @[RA_Mul.scala 47:10:@643.4]
  assign io_matrix_o_3_17 = FA_14_io_cout; // @[RA_Mul.scala 47:10:@659.4]
  assign io_matrix_o_3_18 = FA_16_io_cout; // @[RA_Mul.scala 47:10:@675.4]
  assign io_matrix_o_3_19 = FA_18_io_cout; // @[RA_Mul.scala 47:10:@691.4]
  assign io_matrix_o_3_20 = FA_20_io_cout; // @[RA_Mul.scala 47:10:@707.4]
  assign io_matrix_o_3_21 = HA_3_io_cout; // @[RA_Mul.scala 22:10:@722.4]
  assign io_matrix_o_3_22 = 1'h0; // @[RA_Mul.scala 293:19:@741.4]
  assign io_matrix_o_3_23 = io_matrix_i_4_23; // @[RA_Mul.scala 366:22:@751.4]
  assign io_matrix_o_3_24 = 1'h0; // @[RA_Mul.scala 293:19:@761.4]
  assign io_matrix_o_3_25 = 1'h0; // @[RA_Mul.scala 293:19:@771.4]
  assign io_matrix_o_3_26 = 1'h0; // @[RA_Mul.scala 293:19:@781.4]
  assign io_matrix_o_3_27 = 1'h0; // @[RA_Mul.scala 293:19:@784.4]
  assign io_matrix_o_3_28 = 1'h0; // @[RA_Mul.scala 293:19:@788.4]
  assign io_matrix_o_3_29 = 1'h0; // @[RA_Mul.scala 293:19:@799.4]
  assign io_matrix_o_3_30 = 1'h0; // @[RA_Mul.scala 293:19:@802.4]
  assign io_matrix_o_3_31 = 1'h0; // @[RA_Mul.scala 293:19:@806.4]
  assign HA_io_a = io_matrix_i_0_1; // @[RA_Mul.scala 19:14:@490.4]
  assign HA_io_b = io_matrix_i_1_1; // @[RA_Mul.scala 20:14:@491.4]
  assign FA_io_a = io_matrix_i_0_3; // @[RA_Mul.scala 43:14:@504.4]
  assign FA_io_b = io_matrix_i_1_3; // @[RA_Mul.scala 44:14:@505.4]
  assign FA_io_cin = io_matrix_i_2_3; // @[RA_Mul.scala 45:16:@506.4]
  assign FA_1_io_a = io_matrix_i_0_6; // @[RA_Mul.scala 43:14:@523.4]
  assign FA_1_io_b = io_matrix_i_1_6; // @[RA_Mul.scala 44:14:@524.4]
  assign FA_1_io_cin = io_matrix_i_2_6; // @[RA_Mul.scala 45:16:@525.4]
  assign FA_2_io_a = io_matrix_i_0_7; // @[RA_Mul.scala 43:14:@534.4]
  assign FA_2_io_b = io_matrix_i_1_7; // @[RA_Mul.scala 44:14:@535.4]
  assign FA_2_io_cin = io_matrix_i_2_7; // @[RA_Mul.scala 45:16:@536.4]
  assign FA_3_io_a = io_matrix_i_0_8; // @[RA_Mul.scala 43:14:@544.4]
  assign FA_3_io_b = io_matrix_i_1_8; // @[RA_Mul.scala 44:14:@545.4]
  assign FA_3_io_cin = io_matrix_i_2_8; // @[RA_Mul.scala 45:16:@546.4]
  assign FA_4_io_a = io_matrix_i_0_9; // @[RA_Mul.scala 43:14:@554.4]
  assign FA_4_io_b = io_matrix_i_1_9; // @[RA_Mul.scala 44:14:@555.4]
  assign FA_4_io_cin = io_matrix_i_2_9; // @[RA_Mul.scala 45:16:@556.4]
  assign FA_5_io_a = io_matrix_i_0_10; // @[RA_Mul.scala 43:14:@564.4]
  assign FA_5_io_b = io_matrix_i_1_10; // @[RA_Mul.scala 44:14:@565.4]
  assign FA_5_io_cin = io_matrix_i_2_10; // @[RA_Mul.scala 45:16:@566.4]
  assign FA_6_io_a = io_matrix_i_0_11; // @[RA_Mul.scala 43:14:@574.4]
  assign FA_6_io_b = io_matrix_i_1_11; // @[RA_Mul.scala 44:14:@575.4]
  assign FA_6_io_cin = io_matrix_i_2_11; // @[RA_Mul.scala 45:16:@576.4]
  assign FA_7_io_a = io_matrix_i_0_12; // @[RA_Mul.scala 43:14:@584.4]
  assign FA_7_io_b = io_matrix_i_1_12; // @[RA_Mul.scala 44:14:@585.4]
  assign FA_7_io_cin = io_matrix_i_2_12; // @[RA_Mul.scala 45:16:@586.4]
  assign FA_8_io_a = io_matrix_i_3_12; // @[RA_Mul.scala 43:14:@592.4]
  assign FA_8_io_b = io_matrix_i_4_12; // @[RA_Mul.scala 44:14:@593.4]
  assign FA_8_io_cin = io_matrix_i_5_12; // @[RA_Mul.scala 45:16:@594.4]
  assign FA_9_io_a = io_matrix_i_0_13; // @[RA_Mul.scala 43:14:@601.4]
  assign FA_9_io_b = io_matrix_i_1_13; // @[RA_Mul.scala 44:14:@602.4]
  assign FA_9_io_cin = io_matrix_i_2_13; // @[RA_Mul.scala 45:16:@603.4]
  assign HA_1_io_a = io_matrix_i_3_13; // @[RA_Mul.scala 19:14:@609.4]
  assign HA_1_io_b = io_matrix_i_4_13; // @[RA_Mul.scala 20:14:@610.4]
  assign FA_10_io_a = io_matrix_i_0_14; // @[RA_Mul.scala 43:14:@616.4]
  assign FA_10_io_b = io_matrix_i_1_14; // @[RA_Mul.scala 44:14:@617.4]
  assign FA_10_io_cin = io_matrix_i_2_14; // @[RA_Mul.scala 45:16:@618.4]
  assign HA_2_io_a = io_matrix_i_3_14; // @[RA_Mul.scala 19:14:@624.4]
  assign HA_2_io_b = io_matrix_i_4_14; // @[RA_Mul.scala 20:14:@625.4]
  assign FA_11_io_a = io_matrix_i_0_15; // @[RA_Mul.scala 43:14:@631.4]
  assign FA_11_io_b = io_matrix_i_1_15; // @[RA_Mul.scala 44:14:@632.4]
  assign FA_11_io_cin = io_matrix_i_2_15; // @[RA_Mul.scala 45:16:@633.4]
  assign FA_12_io_a = io_matrix_i_3_15; // @[RA_Mul.scala 43:14:@639.4]
  assign FA_12_io_b = io_matrix_i_4_15; // @[RA_Mul.scala 44:14:@640.4]
  assign FA_12_io_cin = io_matrix_i_5_15; // @[RA_Mul.scala 45:16:@641.4]
  assign FA_13_io_a = io_matrix_i_0_16; // @[RA_Mul.scala 43:14:@647.4]
  assign FA_13_io_b = io_matrix_i_1_16; // @[RA_Mul.scala 44:14:@648.4]
  assign FA_13_io_cin = io_matrix_i_2_16; // @[RA_Mul.scala 45:16:@649.4]
  assign FA_14_io_a = io_matrix_i_3_16; // @[RA_Mul.scala 43:14:@655.4]
  assign FA_14_io_b = io_matrix_i_4_16; // @[RA_Mul.scala 44:14:@656.4]
  assign FA_14_io_cin = io_matrix_i_5_16; // @[RA_Mul.scala 45:16:@657.4]
  assign FA_15_io_a = io_matrix_i_0_17; // @[RA_Mul.scala 43:14:@663.4]
  assign FA_15_io_b = io_matrix_i_1_17; // @[RA_Mul.scala 44:14:@664.4]
  assign FA_15_io_cin = io_matrix_i_2_17; // @[RA_Mul.scala 45:16:@665.4]
  assign FA_16_io_a = io_matrix_i_3_17; // @[RA_Mul.scala 43:14:@671.4]
  assign FA_16_io_b = io_matrix_i_4_17; // @[RA_Mul.scala 44:14:@672.4]
  assign FA_16_io_cin = io_matrix_i_5_17; // @[RA_Mul.scala 45:16:@673.4]
  assign FA_17_io_a = io_matrix_i_0_18; // @[RA_Mul.scala 43:14:@679.4]
  assign FA_17_io_b = io_matrix_i_1_18; // @[RA_Mul.scala 44:14:@680.4]
  assign FA_17_io_cin = io_matrix_i_2_18; // @[RA_Mul.scala 45:16:@681.4]
  assign FA_18_io_a = io_matrix_i_3_18; // @[RA_Mul.scala 43:14:@687.4]
  assign FA_18_io_b = io_matrix_i_4_18; // @[RA_Mul.scala 44:14:@688.4]
  assign FA_18_io_cin = io_matrix_i_5_18; // @[RA_Mul.scala 45:16:@689.4]
  assign FA_19_io_a = io_matrix_i_0_19; // @[RA_Mul.scala 43:14:@695.4]
  assign FA_19_io_b = io_matrix_i_1_19; // @[RA_Mul.scala 44:14:@696.4]
  assign FA_19_io_cin = io_matrix_i_2_19; // @[RA_Mul.scala 45:16:@697.4]
  assign FA_20_io_a = io_matrix_i_3_19; // @[RA_Mul.scala 43:14:@703.4]
  assign FA_20_io_b = io_matrix_i_4_19; // @[RA_Mul.scala 44:14:@704.4]
  assign FA_20_io_cin = io_matrix_i_5_19; // @[RA_Mul.scala 45:16:@705.4]
  assign FA_21_io_a = io_matrix_i_0_20; // @[RA_Mul.scala 43:14:@711.4]
  assign FA_21_io_b = io_matrix_i_1_20; // @[RA_Mul.scala 44:14:@712.4]
  assign FA_21_io_cin = io_matrix_i_2_20; // @[RA_Mul.scala 45:16:@713.4]
  assign HA_3_io_a = io_matrix_i_3_20; // @[RA_Mul.scala 19:14:@719.4]
  assign HA_3_io_b = io_matrix_i_4_20; // @[RA_Mul.scala 20:14:@720.4]
  assign FA_22_io_a = io_matrix_i_0_21; // @[RA_Mul.scala 43:14:@726.4]
  assign FA_22_io_b = io_matrix_i_1_21; // @[RA_Mul.scala 44:14:@727.4]
  assign FA_22_io_cin = io_matrix_i_2_21; // @[RA_Mul.scala 45:16:@728.4]
  assign FA_23_io_a = io_matrix_i_0_22; // @[RA_Mul.scala 43:14:@735.4]
  assign FA_23_io_b = io_matrix_i_1_22; // @[RA_Mul.scala 44:14:@736.4]
  assign FA_23_io_cin = io_matrix_i_2_22; // @[RA_Mul.scala 45:16:@737.4]
  assign FA_24_io_a = io_matrix_i_0_23; // @[RA_Mul.scala 43:14:@745.4]
  assign FA_24_io_b = io_matrix_i_1_23; // @[RA_Mul.scala 44:14:@746.4]
  assign FA_24_io_cin = io_matrix_i_2_23; // @[RA_Mul.scala 45:16:@747.4]
  assign FA_25_io_a = io_matrix_i_0_24; // @[RA_Mul.scala 43:14:@755.4]
  assign FA_25_io_b = io_matrix_i_1_24; // @[RA_Mul.scala 44:14:@756.4]
  assign FA_25_io_cin = io_matrix_i_2_24; // @[RA_Mul.scala 45:16:@757.4]
  assign FA_26_io_a = io_matrix_i_0_25; // @[RA_Mul.scala 43:14:@765.4]
  assign FA_26_io_b = io_matrix_i_1_25; // @[RA_Mul.scala 44:14:@766.4]
  assign FA_26_io_cin = io_matrix_i_2_25; // @[RA_Mul.scala 45:16:@767.4]
  assign FA_27_io_a = io_matrix_i_0_26; // @[RA_Mul.scala 43:14:@775.4]
  assign FA_27_io_b = io_matrix_i_1_26; // @[RA_Mul.scala 44:14:@776.4]
  assign FA_27_io_cin = io_matrix_i_2_26; // @[RA_Mul.scala 45:16:@777.4]
  assign FA_28_io_a = io_matrix_i_0_29; // @[RA_Mul.scala 43:14:@792.4]
  assign FA_28_io_b = io_matrix_i_1_29; // @[RA_Mul.scala 44:14:@793.4]
  assign FA_28_io_cin = io_matrix_i_2_29; // @[RA_Mul.scala 45:16:@794.4]
endmodule
